module boot_rom (
  input          clk,
  input          en,
  input  [11:0]  addr_i,
  output [31:0]  dout_o
);

 // Based on this UG - https://www.xilinx.com/support/documentation/sw_manuals/xilinx2020_1/ug901-vivado-synthesis.pdf

 (*rom_style = "block" *) logic [31:0] data;
 assign dout_o = data;

 always @(posedge clk) begin
     if (en) begin
         case (addr_i)
         'd0: data <= 32'h30005073;         'd1: data <= 32'h70008117;
         'd2: data <= 32'hff810113;         'd3: data <= 32'h70001197;
         'd4: data <= 32'h80c18193;         'd5: data <= 32'h00000517;
         'd6: data <= 32'h12850513;         'd7: data <= 32'h30551073;
         'd8: data <= 32'h30001073;         'd9: data <= 32'h30401073;
         'd10: data <= 32'h00000213;         'd11: data <= 32'h00000293;
         'd12: data <= 32'h00000313;         'd13: data <= 32'h00000393;
         'd14: data <= 32'h00000813;         'd15: data <= 32'h00000893;
         'd16: data <= 32'h00000913;         'd17: data <= 32'h00000993;
         'd18: data <= 32'h00000a13;         'd19: data <= 32'h00000a93;
         'd20: data <= 32'h00000b13;         'd21: data <= 32'h00000b93;
         'd22: data <= 32'h00000c13;         'd23: data <= 32'h00000c93;
         'd24: data <= 32'h00000d13;         'd25: data <= 32'h00000d93;
         'd26: data <= 32'h00000e13;         'd27: data <= 32'h00000e93;
         'd28: data <= 32'h00000f13;         'd29: data <= 32'h00000f93;
         'd30: data <= 32'h00003597;         'd31: data <= 32'h6e058593;
         'd32: data <= 32'h70000617;         'd33: data <= 32'hf8060613;
         'd34: data <= 32'h70000697;         'd35: data <= 32'hf9068693;
         'd36: data <= 32'h00c58e63;         'd37: data <= 32'h00d65c63;
         'd38: data <= 32'h0005a703;         'd39: data <= 32'h00e62023;
         'd40: data <= 32'h00458593;         'd41: data <= 32'h00460613;
         'd42: data <= 32'hfedff06f;         'd43: data <= 32'h70000717;
         'd44: data <= 32'hf7470713;         'd45: data <= 32'h70002797;
         'd46: data <= 32'hf1c78793;         'd47: data <= 32'h00f75863;
         'd48: data <= 32'h00072023;         'd49: data <= 32'h00470713;
         'd50: data <= 32'hff5ff06f;         'd51: data <= 32'h00003417;
         'd52: data <= 32'h32440413;         'd53: data <= 32'h00003497;
         'd54: data <= 32'h31c48493;         'd55: data <= 32'h00945a63;
         'd56: data <= 32'h0009a083;         'd57: data <= 32'h000080e7;
         'd58: data <= 32'h00440413;         'd59: data <= 32'hff1ff06f;
         'd60: data <= 32'h00000513;         'd61: data <= 32'h00000593;
         'd62: data <= 32'h23c000ef;         'd63: data <= 32'h30047073;
         'd64: data <= 32'h34051073;         'd65: data <= 32'h00003417;
         'd66: data <= 32'h2ec40413;         'd67: data <= 32'h00003497;
         'd68: data <= 32'h2e448493;         'd69: data <= 32'h00945a63;
         'd70: data <= 32'h00042083;         'd71: data <= 32'h000080e7;
         'd72: data <= 32'h00440413;         'd73: data <= 32'hff1ff06f;
         'd74: data <= 32'h00000093;         'd75: data <= 32'h00008463;
         'd76: data <= 32'h000080e7;         'd77: data <= 32'h10500073;
         'd78: data <= 32'h0000006f;         'd79: data <= 32'hff810113;
         'd80: data <= 32'h00812023;         'd81: data <= 32'h00912223;
         'd82: data <= 32'h34202473;         'd83: data <= 32'h02044663;
         'd84: data <= 32'h34102473;         'd85: data <= 32'h00041483;
         'd86: data <= 32'h0034f493;         'd87: data <= 32'h00240413;
         'd88: data <= 32'h34141073;         'd89: data <= 32'h00300413;
         'd90: data <= 32'h00941863;         'd91: data <= 32'h34102473;
         'd92: data <= 32'h00240413;         'd93: data <= 32'h34141073;
         'd94: data <= 32'h00012403;         'd95: data <= 32'h00412483;
         'd96: data <= 32'h00810113;         'd97: data <= 32'h30200073;
         'd98: data <= 32'hff010113;         'd99: data <= 32'h00112623;
         'd100: data <= 32'h00812423;         'd101: data <= 32'h00000413;
         'd102: data <= 32'h00040593;         'd103: data <= 32'h00003517;
         'd104: data <= 32'h25450513;         'd105: data <= 32'h4cc000ef;
         'd106: data <= 32'h00a40413;         'd107: data <= 32'h0ff47413;
         'd108: data <= 32'h12c00513;         'd109: data <= 32'h2a0010ef;
         'd110: data <= 32'hfe1ff06f;         'd111: data <= 32'hff010113;
         'd112: data <= 32'h00112623;         'd113: data <= 32'h00812423;
         'd114: data <= 32'h00000413;         'd115: data <= 32'h00040593;
         'd116: data <= 32'h00003517;         'd117: data <= 32'h23850513;
         'd118: data <= 32'h498000ef;         'd119: data <= 32'h00a40413;
         'd120: data <= 32'h0ff47413;         'd121: data <= 32'h09600513;
         'd122: data <= 32'h26c010ef;         'd123: data <= 32'hfe1ff06f;
         'd124: data <= 32'hff010113;         'd125: data <= 32'h00112623;
         'd126: data <= 32'h00812423;         'd127: data <= 32'h00000413;
         'd128: data <= 32'h00040593;         'd129: data <= 32'h00003517;
         'd130: data <= 32'h21c50513;         'd131: data <= 32'h464000ef;
         'd132: data <= 32'h00440413;         'd133: data <= 32'h0ff47413;
         'd134: data <= 32'h06400513;         'd135: data <= 32'h238010ef;
         'd136: data <= 32'hfe1ff06f;         'd137: data <= 32'hff010113;
         'd138: data <= 32'h00112623;         'd139: data <= 32'h00812423;
         'd140: data <= 32'h00000413;         'd141: data <= 32'h00040593;
         'd142: data <= 32'h00003517;         'd143: data <= 32'h20050513;
         'd144: data <= 32'h430000ef;         'd145: data <= 32'h00240413;
         'd146: data <= 32'h0ff47413;         'd147: data <= 32'h03200513;
         'd148: data <= 32'h204010ef;         'd149: data <= 32'hfe1ff06f;
         'd150: data <= 32'hfe010113;         'd151: data <= 32'h00112e23;
         'd152: data <= 32'h00012623;         'd153: data <= 32'h00012423;
         'd154: data <= 32'h00012223;         'd155: data <= 32'h00012023;
         'd156: data <= 32'h00c10793;         'd157: data <= 32'h00100713;
         'd158: data <= 32'h00000693;         'd159: data <= 32'h10000613;
         'd160: data <= 32'h00003597;         'd161: data <= 32'h1d058593;
         'd162: data <= 32'h00000517;         'd163: data <= 32'hf9c50513;
         'd164: data <= 32'h345000ef;         'd165: data <= 32'h00810793;
         'd166: data <= 32'h00100713;         'd167: data <= 32'h00000693;
         'd168: data <= 32'h10000613;         'd169: data <= 32'h00003597;
         'd170: data <= 32'h1b058593;         'd171: data <= 32'h00000517;
         'd172: data <= 32'hf4450513;         'd173: data <= 32'h321000ef;
         'd174: data <= 32'h00410793;         'd175: data <= 32'h00100713;
         'd176: data <= 32'h00000693;         'd177: data <= 32'h10000613;
         'd178: data <= 32'h00003597;         'd179: data <= 32'h19058593;
         'd180: data <= 32'h00000517;         'd181: data <= 32'heec50513;
         'd182: data <= 32'h2fd000ef;         'd183: data <= 32'h00010793;
         'd184: data <= 32'h00100713;         'd185: data <= 32'h00000693;
         'd186: data <= 32'h10000613;         'd187: data <= 32'h00003597;
         'd188: data <= 32'h17058593;         'd189: data <= 32'h00000517;
         'd190: data <= 32'he9450513;         'd191: data <= 32'h2d9000ef;
         'd192: data <= 32'h3b9000ef;         'd193: data <= 32'h0000006f;
         'd194: data <= 32'hff010113;         'd195: data <= 32'h00112623;
         'd196: data <= 32'h00003797;         'd197: data <= 32'hef078793;
         'd198: data <= 32'h30579073;         'd199: data <= 32'h0001c537;
         'd200: data <= 32'h20050513;         'd201: data <= 32'h284000ef;
         'd202: data <= 32'h00c12083;         'd203: data <= 32'h01010113;
         'd204: data <= 32'h00008067;         'd205: data <= 32'hff010113;
         'd206: data <= 32'h00112623;         'd207: data <= 32'hfcdff0ef;
         'd208: data <= 32'h00003597;         'd209: data <= 32'h12058593;
         'd210: data <= 32'h00003517;         'd211: data <= 32'h12450513;
         'd212: data <= 32'h320000ef;         'd213: data <= 32'hf05ff0ef;
         'd214: data <= 32'h00c12083;         'd215: data <= 32'h01010113;
         'd216: data <= 32'h00008067;         'd217: data <= 32'hff010113;
         'd218: data <= 32'h00112623;         'd219: data <= 32'h34405073;
         'd220: data <= 32'h34405073;         'd221: data <= 32'h34405073;
         'd222: data <= 32'h28c000ef;         'd223: data <= 32'h00050593;
         'd224: data <= 32'h00003517;         'd225: data <= 32'h10c50513;
         'd226: data <= 32'h2e8000ef;         'd227: data <= 32'h342025f3;
         'd228: data <= 32'h00003517;         'd229: data <= 32'h10450513;
         'd230: data <= 32'h2d8000ef;         'd231: data <= 32'h00c12083;
         'd232: data <= 32'h01010113;         'd233: data <= 32'h00008067;
         'd234: data <= 32'hff010113;         'd235: data <= 32'h00112623;
         'd236: data <= 32'h342025f3;         'd237: data <= 32'h00003517;
         'd238: data <= 32'h10050513;         'd239: data <= 32'h2b4000ef;
         'd240: data <= 32'h00c12083;         'd241: data <= 32'h01010113;
         'd242: data <= 32'h00008067;         'd243: data <= 32'hff010113;
         'd244: data <= 32'h00112623;         'd245: data <= 32'h30047073;
         'd246: data <= 32'h00003517;         'd247: data <= 32'h0fc50513;
         'd248: data <= 32'h23c000ef;         'd249: data <= 32'h00100073;
         'd250: data <= 32'h0000006f;         'd251: data <= 32'h00008067;
         'd252: data <= 32'hff010113;         'd253: data <= 32'h00112623;
         'd254: data <= 32'h30047073;         'd255: data <= 32'h00003517;
         'd256: data <= 32'h14850513;         'd257: data <= 32'h218000ef;
         'd258: data <= 32'h00100073;         'd259: data <= 32'h0000006f;
         'd260: data <= 32'h00008067;         'd261: data <= 32'hfe010113;
         'd262: data <= 32'h00112e23;         'd263: data <= 32'h00812c23;
         'd264: data <= 32'h00912a23;         'd265: data <= 32'h01212823;
         'd266: data <= 32'h00050493;         'd267: data <= 32'h00058913;
         'd268: data <= 32'h00010723;         'd269: data <= 32'h00058523;
         'd270: data <= 32'h00000413;         'd271: data <= 32'h0480006f;
         'd272: data <= 32'h00a00593;         'd273: data <= 32'h00048513;
         'd274: data <= 32'h2e5020ef;         'd275: data <= 32'h00003797;
         'd276: data <= 32'h1c078793;         'd277: data <= 32'h00a787b3;
         'd278: data <= 32'h0007c703;         'd279: data <= 32'h01040793;
         'd280: data <= 32'h002787b3;         'd281: data <= 32'hfee78a23;
         'd282: data <= 32'h00a00593;         'd283: data <= 32'h00048513;
         'd284: data <= 32'h275020ef;         'd285: data <= 32'h00050493;
         'd286: data <= 32'h00140413;         'd287: data <= 32'h01041413;
         'd288: data <= 32'h01045413;         'd289: data <= 32'h00900793;
         'd290: data <= 32'hfa87fce3;         'd291: data <= 32'h02078a63;
         'd292: data <= 32'h01078713;         'd293: data <= 32'h00270733;
         'd294: data <= 32'hff474683;         'd295: data <= 32'h03000713;
         'd296: data <= 32'h02e69463;         'd297: data <= 32'h01078713;
         'd298: data <= 32'h00270733;         'd299: data <= 32'hfe070a23;
         'd300: data <= 32'hfff78793;         'd301: data <= 32'h01079793;
         'd302: data <= 32'h0107d793;         'd303: data <= 32'hfd1ff06f;
         'd304: data <= 32'h00078693;         'd305: data <= 32'h0200006f;
         'd306: data <= 32'h00000693;         'd307: data <= 32'h0180006f;
         'd308: data <= 32'hfff78713;         'd309: data <= 32'h01071713;
         'd310: data <= 32'h01075713;         'd311: data <= 32'h02078863;
         'd312: data <= 32'h00070793;         'd313: data <= 32'h01078713;
         'd314: data <= 32'h00270733;         'd315: data <= 32'hff474703;
         'd316: data <= 32'hfe0700e3;         'd317: data <= 32'h00168613;
         'd318: data <= 32'h00d906b3;         'd319: data <= 32'h00e68023;
         'd320: data <= 32'h01061693;         'd321: data <= 32'h0106d693;
         'd322: data <= 32'hfc9ff06f;         'd323: data <= 32'h00d90933;
         'd324: data <= 32'h00090023;         'd325: data <= 32'h01c12083;
         'd326: data <= 32'h01812403;         'd327: data <= 32'h01412483;
         'd328: data <= 32'h01012903;         'd329: data <= 32'h02010113;
         'd330: data <= 32'h00008067;         'd331: data <= 32'h00000693;
         'd332: data <= 32'h0340006f;         'd333: data <= 32'h00269713;
         'd334: data <= 32'h00e55733;         'd335: data <= 32'h00f77713;
         'd336: data <= 32'h00700793;         'd337: data <= 32'h40d787b3;
         'd338: data <= 32'h00f587b3;         'd339: data <= 32'h00003617;
         'd340: data <= 32'h0ac60613;         'd341: data <= 32'h00e60733;
         'd342: data <= 32'h00074703;         'd343: data <= 32'h00e78023;
         'd344: data <= 32'h00168693;         'd345: data <= 32'h00700793;
         'd346: data <= 32'hfcd7d6e3;         'd347: data <= 32'h00058423;
         'd348: data <= 32'h00008067;         'd349: data <= 32'h00c0006f;
         'd350: data <= 32'h00158593;         'd351: data <= 32'hfff50513;
         'd352: data <= 32'h02050263;         'd353: data <= 32'h0005c703;
         'd354: data <= 32'hf9f70793;         'd355: data <= 32'h0ff7f793;
         'd356: data <= 32'h01900693;         'd357: data <= 32'hfef6e2e3;
         'd358: data <= 32'hfe070713;         'd359: data <= 32'h00e58023;
         'd360: data <= 32'hfd9ff06f;         'd361: data <= 32'h00008067;
         'd362: data <= 32'hff010113;         'd363: data <= 32'h00112623;
         'd364: data <= 32'h00050593;         'd365: data <= 32'h02faf537;
         'd366: data <= 32'h08050513;         'd367: data <= 32'h129020ef;
         'd368: data <= 32'hb00007b7;         'd369: data <= 32'h00a7a023;
         'd370: data <= 32'h00c12083;         'd371: data <= 32'h01010113;
         'd372: data <= 32'h00008067;         'd373: data <= 32'hb00007b7;
         'd374: data <= 32'h0047a783;         'd375: data <= 32'h00010737;
         'd376: data <= 32'h00e7f7b3;         'd377: data <= 32'hfe0788e3;
         'd378: data <= 32'hb00007b7;         'd379: data <= 32'h00a7a623;
         'd380: data <= 32'h00008067;         'd381: data <= 32'hb00007b7;
         'd382: data <= 32'h0087a503;         'd383: data <= 32'h0ff57513;
         'd384: data <= 32'h00008067;         'd385: data <= 32'hff010113;
         'd386: data <= 32'h00112623;         'd387: data <= 32'hfe9ff0ef;
         'd388: data <= 32'h00c12083;         'd389: data <= 32'h01010113;
         'd390: data <= 32'h00008067;         'd391: data <= 32'hff010113;
         'd392: data <= 32'h00112623;         'd393: data <= 32'h00812423;
         'd394: data <= 32'h00912223;         'd395: data <= 32'h0100006f;
         'd396: data <= 32'h00040513;         'd397: data <= 32'hfa1ff0ef;
         'd398: data <= 32'h00048513;         'd399: data <= 32'h00150493;
         'd400: data <= 32'h00054403;         'd401: data <= 32'h00040c63;
         'd402: data <= 32'h00a00793;         'd403: data <= 32'hfef412e3;
         'd404: data <= 32'h00d00513;         'd405: data <= 32'hf81ff0ef;
         'd406: data <= 32'hfd9ff06f;         'd407: data <= 32'h00c12083;
         'd408: data <= 32'h00812403;         'd409: data <= 32'h00412483;
         'd410: data <= 32'h01010113;         'd411: data <= 32'h00008067;
         'd412: data <= 32'hfc010113;         'd413: data <= 32'h00112e23;
         'd414: data <= 32'h00812c23;         'd415: data <= 32'h00912a23;
         'd416: data <= 32'h01212823;         'd417: data <= 32'h00050493;
         'd418: data <= 32'h02b12223;         'd419: data <= 32'h02c12423;
         'd420: data <= 32'h02d12623;         'd421: data <= 32'h02e12823;
         'd422: data <= 32'h02f12a23;         'd423: data <= 32'h03012c23;
         'd424: data <= 32'h03112e23;         'd425: data <= 32'h02410793;
         'd426: data <= 32'h00f12023;         'd427: data <= 32'h1240006f;
         'd428: data <= 32'h00248493;         'd429: data <= 32'h00094403;
         'd430: data <= 32'hfa840793;         'd431: data <= 32'h0ff7f693;
         'd432: data <= 32'h02000713;         'd433: data <= 32'h0ed76663;
         'd434: data <= 32'h00269793;         'd435: data <= 32'h00003717;
         'd436: data <= 32'hea870713;         'd437: data <= 32'h00e787b3;
         'd438: data <= 32'h0007a783;         'd439: data <= 32'h00e787b3;
         'd440: data <= 32'h00078067;         'd441: data <= 32'h00012783;
         'd442: data <= 32'h00478713;         'd443: data <= 32'h00e12023;
         'd444: data <= 32'h0007a503;         'd445: data <= 32'hf29ff0ef;
         'd446: data <= 32'h0d80006f;         'd447: data <= 32'h00012783;
         'd448: data <= 32'h00478713;         'd449: data <= 32'h00e12023;
         'd450: data <= 32'h0007c503;         'd451: data <= 32'hec9ff0ef;
         'd452: data <= 32'h0c00006f;         'd453: data <= 32'h00012783;
         'd454: data <= 32'h00478713;         'd455: data <= 32'h00e12023;
         'd456: data <= 32'h0007a403;         'd457: data <= 32'h00044e63;
         'd458: data <= 32'h00410593;         'd459: data <= 32'h00040513;
         'd460: data <= 32'hce5ff0ef;         'd461: data <= 32'h00410513;
         'd462: data <= 32'hee5ff0ef;         'd463: data <= 32'h0940006f;
         'd464: data <= 32'h40800433;         'd465: data <= 32'h02d00513;
         'd466: data <= 32'he8dff0ef;         'd467: data <= 32'hfddff06f;
         'd468: data <= 32'h00012783;         'd469: data <= 32'h00478713;
         'd470: data <= 32'h00e12023;         'd471: data <= 32'h00410593;
         'd472: data <= 32'h0007a503;         'd473: data <= 32'hcb1ff0ef;
         'd474: data <= 32'h00410513;         'd475: data <= 32'heb1ff0ef;
         'd476: data <= 32'h0600006f;         'd477: data <= 32'h00012783;
         'd478: data <= 32'h00478713;         'd479: data <= 32'h00e12023;
         'd480: data <= 32'h00410593;         'd481: data <= 32'h0007a503;
         'd482: data <= 32'hda5ff0ef;         'd483: data <= 32'h05800793;
         'd484: data <= 32'h00f40863;         'd485: data <= 32'h00410513;
         'd486: data <= 32'he85ff0ef;         'd487: data <= 32'h0340006f;
         'd488: data <= 32'h00410593;         'd489: data <= 32'h00b00513;
         'd490: data <= 32'hdcdff0ef;         'd491: data <= 32'hfe9ff06f;
         'd492: data <= 32'h02500513;         'd493: data <= 32'he21ff0ef;
         'd494: data <= 32'h00040513;         'd495: data <= 32'he19ff0ef;
         'd496: data <= 32'h0100006f;         'd497: data <= 32'h00040513;
         'd498: data <= 32'he0dff0ef;         'd499: data <= 32'h00090493;
         'd500: data <= 32'h00148913;         'd501: data <= 32'h0004c403;
         'd502: data <= 32'h02040063;         'd503: data <= 32'h02500793;
         'd504: data <= 32'hecf408e3;         'd505: data <= 32'h00a00793;
         'd506: data <= 32'hfcf41ee3;         'd507: data <= 32'h00d00513;
         'd508: data <= 32'hde5ff0ef;         'd509: data <= 32'hfd1ff06f;
         'd510: data <= 32'h01c12083;         'd511: data <= 32'h01812403;
         'd512: data <= 32'h01412483;         'd513: data <= 32'h01012903;
         'd514: data <= 32'h04010113;         'd515: data <= 32'h00008067;
         'd516: data <= 32'h70000797;         'd517: data <= 32'h8447a783;
         'd518: data <= 32'h0007a783;         'd519: data <= 32'h00079a63;
         'd520: data <= 32'hfff00793;         'd521: data <= 32'h70000717;
         'd522: data <= 32'h80f72223;         'd523: data <= 32'h00008067;
         'd524: data <= 32'h70000797;         'd525: data <= 32'h8247a783;
         'd526: data <= 32'h00c7a783;         'd527: data <= 32'h0007a783;
         'd528: data <= 32'h6ffff717;         'd529: data <= 32'h7ef72423;
         'd530: data <= 32'h00008067;         'd531: data <= 32'hff010113;
         'd532: data <= 32'h00112623;         'd533: data <= 32'h00812423;
         'd534: data <= 32'h00050413;         'd535: data <= 32'h03052503;
         'd536: data <= 32'h1f9010ef;         'd537: data <= 32'h00040513;
         'd538: data <= 32'h1f1010ef;         'd539: data <= 32'h00c12083;
         'd540: data <= 32'h00812403;         'd541: data <= 32'h01010113;
         'd542: data <= 32'h00008067;         'd543: data <= 32'hfe010113;
         'd544: data <= 32'h00112e23;         'd545: data <= 32'h00812c23;
         'd546: data <= 32'h00912a23;         'd547: data <= 32'h01212823;
         'd548: data <= 32'h01312623;         'd549: data <= 32'h01412423;
         'd550: data <= 32'h01512223;         'd551: data <= 32'h01612023;
         'd552: data <= 32'h00050a93;         'd553: data <= 32'h00058493;
         'd554: data <= 32'h00060913;         'd555: data <= 32'h00068b13;
         'd556: data <= 32'h00070993;         'd557: data <= 32'h00078a13;
         'd558: data <= 32'h00080413;         'd559: data <= 32'h00261613;
         'd560: data <= 32'h0a500593;         'd561: data <= 32'h03082503;
         'd562: data <= 32'h4c8020ef;         'd563: data <= 32'h03042703;
         'd564: data <= 32'h400007b7;         'd565: data <= 32'hfff78793;
         'd566: data <= 32'h00f907b3;         'd567: data <= 32'h00279793;
         'd568: data <= 32'h00f707b3;         'd569: data <= 32'hff07f913;
         'd570: data <= 32'h02048863;         'd571: data <= 32'h00000613;
         'd572: data <= 32'h00f00813;         'd573: data <= 32'h02c86063;
         'd574: data <= 32'h00c48833;         'd575: data <= 32'h00084883;
         'd576: data <= 32'h00c40833;         'd577: data <= 32'h03180a23;
         'd578: data <= 32'h00088663;         'd579: data <= 32'h00160613;
         'd580: data <= 32'hfe1ff06f;         'd581: data <= 32'h040401a3;
         'd582: data <= 32'h00400793;         'd583: data <= 32'h0137f863;
         'd584: data <= 32'h30047073;         'd585: data <= 32'h00100073;
         'd586: data <= 32'h0000006f;         'd587: data <= 32'h03342623;
         'd588: data <= 32'h05342223;         'd589: data <= 32'h00440513;
         'd590: data <= 32'h1f1010ef;         'd591: data <= 32'h01840513;
         'd592: data <= 32'h1e9010ef;         'd593: data <= 32'h00842823;
         'd594: data <= 32'h00500793;         'd595: data <= 32'h413787b3;
         'd596: data <= 32'h00f42c23;         'd597: data <= 32'h02842223;
         'd598: data <= 32'h000b0613;         'd599: data <= 32'h000a8593;
         'd600: data <= 32'h00090513;         'd601: data <= 32'h70c020ef;
         'd602: data <= 32'h00a42023;         'd603: data <= 32'h000a0463;
         'd604: data <= 32'h008a2023;         'd605: data <= 32'h01c12083;
         'd606: data <= 32'h01812403;         'd607: data <= 32'h01412483;
         'd608: data <= 32'h01012903;         'd609: data <= 32'h00c12983;
         'd610: data <= 32'h00812a03;         'd611: data <= 32'h00412a83;
         'd612: data <= 32'h00012b03;         'd613: data <= 32'h02010113;
         'd614: data <= 32'h00008067;         'd615: data <= 32'hff010113;
         'd616: data <= 32'h00112623;         'd617: data <= 32'h00812423;
         'd618: data <= 32'h00000413;         'd619: data <= 32'h0240006f;
         'd620: data <= 32'h00241793;         'd621: data <= 32'h008787b3;
         'd622: data <= 32'h00279713;         'd623: data <= 32'h6ffff517;
         'd624: data <= 32'h74850513;         'd625: data <= 32'h00e50533;
         'd626: data <= 32'h141010ef;         'd627: data <= 32'h00140413;
         'd628: data <= 32'h00400793;         'd629: data <= 32'hfc87fee3;
         'd630: data <= 32'h6ffff517;         'd631: data <= 32'h71850513;
         'd632: data <= 32'h129010ef;         'd633: data <= 32'h6ffff517;
         'd634: data <= 32'h6f850513;         'd635: data <= 32'h11d010ef;
         'd636: data <= 32'h6ffff517;         'd637: data <= 32'h6d850513;
         'd638: data <= 32'h111010ef;         'd639: data <= 32'h6ffff517;
         'd640: data <= 32'h6b850513;         'd641: data <= 32'h105010ef;
         'd642: data <= 32'h6ffff517;         'd643: data <= 32'h69850513;
         'd644: data <= 32'h0f9010ef;         'd645: data <= 32'h6ffff797;
         'd646: data <= 32'h6dc78793;         'd647: data <= 32'h6ffff717;
         'd648: data <= 32'h62f72c23;         'd649: data <= 32'h6ffff797;
         'd650: data <= 32'h6b878793;         'd651: data <= 32'h6ffff717;
         'd652: data <= 32'h62f72223;         'd653: data <= 32'h00c12083;
         'd654: data <= 32'h00812403;         'd655: data <= 32'h01010113;
         'd656: data <= 32'h00008067;         'd657: data <= 32'hff010113;
         'd658: data <= 32'h00112623;         'd659: data <= 32'h00812423;
         'd660: data <= 32'h00050413;         'd661: data <= 32'h30047073;
         'd662: data <= 32'h6ffff717;         'd663: data <= 32'h5b870713;
         'd664: data <= 32'h00072783;         'd665: data <= 32'h00178793;
         'd666: data <= 32'h00f72023;         'd667: data <= 32'h6ffff717;
         'd668: data <= 32'h5dc70713;         'd669: data <= 32'h00072783;
         'd670: data <= 32'h00178793;         'd671: data <= 32'h00f72023;
         'd672: data <= 32'h6ffff797;         'd673: data <= 32'h5d87a783;
         'd674: data <= 32'h02078863;         'd675: data <= 32'h6ffff797;
         'd676: data <= 32'h5b07a783;         'd677: data <= 32'h02079e63;
         'd678: data <= 32'h6ffff797;         'd679: data <= 32'h5c07a783;
         'd680: data <= 32'h02c7a703;         'd681: data <= 32'h02c52783;
         'd682: data <= 32'h02e7e463;         'd683: data <= 32'h6ffff797;
         'd684: data <= 32'h5aa7a623;         'd685: data <= 32'h01c0006f;
         'd686: data <= 32'h6ffff797;         'd687: data <= 32'h5aa7a023;
         'd688: data <= 32'h6ffff717;         'd689: data <= 32'h58872703;
         'd690: data <= 32'h00100793;         'd691: data <= 32'h0ef70663;
         'd692: data <= 32'h6ffff717;         'd693: data <= 32'h55c70713;
         'd694: data <= 32'h00072783;         'd695: data <= 32'h00178793;
         'd696: data <= 32'h00f72023;         'd697: data <= 32'h02c42703;
         'd698: data <= 32'h00100793;         'd699: data <= 32'h00e797b3;
         'd700: data <= 32'h6ffff697;         'd701: data <= 32'h55068693;
         'd702: data <= 32'h0006a603;         'd703: data <= 32'h00c7e7b3;
         'd704: data <= 32'h00f6a023;         'd705: data <= 32'h6ffff697;
         'd706: data <= 32'h60068693;         'd707: data <= 32'h00271793;
         'd708: data <= 32'h00e787b3;         'd709: data <= 32'h00279793;
         'd710: data <= 32'h00f687b3;         'd711: data <= 32'h0047a783;
         'd712: data <= 32'h00f42423;         'd713: data <= 32'h0087a603;
         'd714: data <= 32'h00c42623;         'd715: data <= 32'h00440713;
         'd716: data <= 32'h00e62223;         'd717: data <= 32'h00e7a423;
         'd718: data <= 32'h02c42603;         'd719: data <= 32'h00261793;
         'd720: data <= 32'h00c78733;         'd721: data <= 32'h00271713;
         'd722: data <= 32'h00d70733;         'd723: data <= 32'h00e42a23;
         'd724: data <= 32'h00072703;         'd725: data <= 32'h00170713;
         'd726: data <= 32'h00c787b3;         'd727: data <= 32'h00279793;
         'd728: data <= 32'h00f686b3;         'd729: data <= 32'h00e6a023;
         'd730: data <= 32'h6ffff717;         'd731: data <= 32'h4a870713;
         'd732: data <= 32'h00072783;         'd733: data <= 32'hfff78793;
         'd734: data <= 32'h00f72023;         'd735: data <= 32'h00079463;
         'd736: data <= 32'h30046073;         'd737: data <= 32'h6ffff797;
         'd738: data <= 32'h4b87a783;         'd739: data <= 32'h00078e63;
         'd740: data <= 32'h6ffff797;         'd741: data <= 32'h4c87a783;
         'd742: data <= 32'h02c7a703;         'd743: data <= 32'h02c42783;
         'd744: data <= 32'h00f77463;         'd745: data <= 32'h00000073;
         'd746: data <= 32'h00c12083;         'd747: data <= 32'h00812403;
         'd748: data <= 32'h01010113;         'd749: data <= 32'h00008067;
         'd750: data <= 32'hde5ff0ef;         'd751: data <= 32'hf15ff06f;
         'd752: data <= 32'h6ffff797;         'd753: data <= 32'h48c7a783;
         'd754: data <= 32'h0a078663;         'd755: data <= 32'hff010113;
         'd756: data <= 32'h00112623;         'd757: data <= 32'h00812423;
         'd758: data <= 32'h00912223;         'd759: data <= 32'h0180006f;
         'd760: data <= 32'h00048513;         'd761: data <= 32'hc69ff0ef;
         'd762: data <= 32'h6ffff797;         'd763: data <= 32'h4647a783;
         'd764: data <= 32'h06078863;         'd765: data <= 32'h30047073;
         'd766: data <= 32'h6ffff417;         'd767: data <= 32'h41840413;
         'd768: data <= 32'h00042783;         'd769: data <= 32'h00178793;
         'd770: data <= 32'h00f42023;         'd771: data <= 32'h6ffff797;
         'd772: data <= 32'h4b47a783;         'd773: data <= 32'h00c7a483;
         'd774: data <= 32'h00448513;         'd775: data <= 32'h764010ef;
         'd776: data <= 32'h6ffff717;         'd777: data <= 32'h42870713;
         'd778: data <= 32'h00072783;         'd779: data <= 32'hfff78793;
         'd780: data <= 32'h00f72023;         'd781: data <= 32'h6ffff717;
         'd782: data <= 32'h41870713;         'd783: data <= 32'h00072783;
         'd784: data <= 32'hfff78793;         'd785: data <= 32'h00f72023;
         'd786: data <= 32'h00042783;         'd787: data <= 32'hfff78793;
         'd788: data <= 32'h00f42023;         'd789: data <= 32'hf80796e3;
         'd790: data <= 32'h30046073;         'd791: data <= 32'hf85ff06f;
         'd792: data <= 32'h00c12083;         'd793: data <= 32'h00812403;
         'd794: data <= 32'h00412483;         'd795: data <= 32'h01010113;
         'd796: data <= 32'h00008067;         'd797: data <= 32'h00008067;
         'd798: data <= 32'hff010113;         'd799: data <= 32'h00112623;
         'd800: data <= 32'h00812423;         'd801: data <= 32'h00912223;
         'd802: data <= 32'h01212023;         'd803: data <= 32'h00050413;
         'd804: data <= 32'h00058493;         'd805: data <= 32'h6ffff917;
         'd806: data <= 32'h3b092903;         'd807: data <= 32'h6ffff797;
         'd808: data <= 32'h3bc78793;         'd809: data <= 32'h0007a703;
         'd810: data <= 32'h06070023;         'd811: data <= 32'h0007a503;
         'd812: data <= 32'h00450513;         'd813: data <= 32'h6cc010ef;
         'd814: data <= 32'h02051863;         'd815: data <= 32'h6ffff797;
         'd816: data <= 32'h39c7a783;         'd817: data <= 32'h02c7a703;
         'd818: data <= 32'h00100793;         'd819: data <= 32'h00e797b3;
         'd820: data <= 32'hfff7c793;         'd821: data <= 32'h6ffff697;
         'd822: data <= 32'h36c68693;         'd823: data <= 32'h0006a703;
         'd824: data <= 32'h00f777b3;         'd825: data <= 32'h00f6a023;
         'd826: data <= 32'hfff00793;         'd827: data <= 32'h04f40463;
         'd828: data <= 32'h00890433;         'd829: data <= 32'h6ffff797;
         'd830: data <= 32'h3647a783;         'd831: data <= 32'h0087a223;
         'd832: data <= 32'h09247863;         'd833: data <= 32'h6ffff517;
         'd834: data <= 32'h34c52503;         'd835: data <= 32'h6ffff597;
         'd836: data <= 32'h34c5a583;         'd837: data <= 32'h00458593;
         'd838: data <= 32'h618010ef;         'd839: data <= 32'h00c12083;
         'd840: data <= 32'h00812403;         'd841: data <= 32'h00412483;
         'd842: data <= 32'h00012903;         'd843: data <= 32'h01010113;
         'd844: data <= 32'h00008067;         'd845: data <= 32'hfa048ee3;
         'd846: data <= 32'h6ffff717;         'd847: data <= 32'h36870713;
         'd848: data <= 32'h00472683;         'd849: data <= 32'h6ffff797;
         'd850: data <= 32'h31478793;         'd851: data <= 32'h0007a603;
         'd852: data <= 32'h00d62423;         'd853: data <= 32'h0007a603;
         'd854: data <= 32'h0086a583;         'd855: data <= 32'h00b62623;
         'd856: data <= 32'h0007a603;         'd857: data <= 32'h00460613;
         'd858: data <= 32'h00c5a223;         'd859: data <= 32'h0007a603;
         'd860: data <= 32'h00460613;         'd861: data <= 32'h00c6a423;
         'd862: data <= 32'h0007a783;         'd863: data <= 32'h00e7aa23;
         'd864: data <= 32'h00072783;         'd865: data <= 32'h00178793;
         'd866: data <= 32'h00f72023;         'd867: data <= 32'hf91ff06f;
         'd868: data <= 32'h6ffff517;         'd869: data <= 32'h2c452503;
         'd870: data <= 32'h6ffff597;         'd871: data <= 32'h2c05a583;
         'd872: data <= 32'h00458593;         'd873: data <= 32'h58c010ef;
         'd874: data <= 32'h6ffff797;         'd875: data <= 32'h2807a783;
         'd876: data <= 32'hf6f476e3;         'd877: data <= 32'h6ffff797;
         'd878: data <= 32'h2687aa23;         'd879: data <= 32'hf61ff06f;
         'd880: data <= 32'hff010113;         'd881: data <= 32'h00112623;
         'd882: data <= 32'hdf9ff0ef;         'd883: data <= 32'he20ff0ef;
         'd884: data <= 32'hff9ff06f;         'd885: data <= 32'hfd010113;
         'd886: data <= 32'h02112623;         'd887: data <= 32'h02812423;
         'd888: data <= 32'h02912223;         'd889: data <= 32'h03212023;
         'd890: data <= 32'h01312e23;         'd891: data <= 32'h01412c23;
         'd892: data <= 32'h01512a23;         'd893: data <= 32'h01612823;
         'd894: data <= 32'h01712623;         'd895: data <= 32'h00050993;
         'd896: data <= 32'h00058a13;         'd897: data <= 32'h00060493;
         'd898: data <= 32'h00068a93;         'd899: data <= 32'h00070b13;
         'd900: data <= 32'h00078b93;         'd901: data <= 32'h00261513;
         'd902: data <= 32'h2a8010ef;         'd903: data <= 32'h06050663;
         'd904: data <= 32'h00050413;         'd905: data <= 32'h06400513;
         'd906: data <= 32'h298010ef;         'd907: data <= 32'h00050913;
         'd908: data <= 32'h04050463;         'd909: data <= 32'h06400613;
         'd910: data <= 32'h00000593;         'd911: data <= 32'h755010ef;
         'd912: data <= 32'h02892823;         'd913: data <= 32'h00000893;
         'd914: data <= 32'h00090813;         'd915: data <= 32'h000b8793;
         'd916: data <= 32'h000b0713;         'd917: data <= 32'h000a8693;
         'd918: data <= 32'h00048613;         'd919: data <= 32'h000a0593;
         'd920: data <= 32'h00098513;         'd921: data <= 32'ha19ff0ef;
         'd922: data <= 32'h00090513;         'd923: data <= 32'hbd9ff0ef;
         'd924: data <= 32'h00100513;         'd925: data <= 32'h0180006f;
         'd926: data <= 32'h00040513;         'd927: data <= 32'h3dc010ef;
         'd928: data <= 32'hfff00513;         'd929: data <= 32'h0080006f;
         'd930: data <= 32'hfff00513;         'd931: data <= 32'h02c12083;
         'd932: data <= 32'h02812403;         'd933: data <= 32'h02412483;
         'd934: data <= 32'h02012903;         'd935: data <= 32'h01c12983;
         'd936: data <= 32'h01812a03;         'd937: data <= 32'h01412a83;
         'd938: data <= 32'h01012b03;         'd939: data <= 32'h00c12b83;
         'd940: data <= 32'h03010113;         'd941: data <= 32'h00008067;
         'd942: data <= 32'hff010113;         'd943: data <= 32'h00112623;
         'd944: data <= 32'h6ffff797;         'd945: data <= 32'h16478793;
         'd946: data <= 32'h00000713;         'd947: data <= 32'h00000693;
         'd948: data <= 32'h08000613;         'd949: data <= 32'h00002597;
         'd950: data <= 32'h74458593;         'd951: data <= 32'h00000517;
         'd952: data <= 32'hee450513;         'd953: data <= 32'hef1ff0ef;
         'd954: data <= 32'h00100793;         'd955: data <= 32'h02f50063;
         'd956: data <= 32'hfff00793;         'd957: data <= 32'h04f50863;
         'd958: data <= 32'h6ffff797;         'd959: data <= 32'h1107a783;
         'd960: data <= 32'h00c12083;         'd961: data <= 32'h01010113;
         'd962: data <= 32'h00008067;         'd963: data <= 32'h050010ef;
         'd964: data <= 32'h00100793;         'd965: data <= 32'hfcf51ee3;
         'd966: data <= 32'h30047073;         'd967: data <= 32'hfff00793;
         'd968: data <= 32'h6ffff717;         'd969: data <= 32'h10f72423;
         'd970: data <= 32'h00100793;         'd971: data <= 32'h6ffff717;
         'd972: data <= 32'h10f72823;         'd973: data <= 32'h6ffff797;
         'd974: data <= 32'h1007a823;         'd975: data <= 32'h0f4020ef;
         'd976: data <= 32'hfb9ff06f;         'd977: data <= 32'h30047073;
         'd978: data <= 32'h00100073;         'd979: data <= 32'h0000006f;
         'd980: data <= 32'h6ffff717;         'd981: data <= 32'h0d070713;
         'd982: data <= 32'h00072783;         'd983: data <= 32'h00178793;
         'd984: data <= 32'h00f72023;         'd985: data <= 32'h00008067;
         'd986: data <= 32'h6ffff517;         'd987: data <= 32'h0dc52503;
         'd988: data <= 32'h00008067;         'd989: data <= 32'hff010113;
         'd990: data <= 32'h00112623;         'd991: data <= 32'h00812423;
         'd992: data <= 32'h00912223;         'd993: data <= 32'h6ffff797;
         'd994: data <= 32'h09c7a783;         'd995: data <= 32'h24079063;
         'd996: data <= 32'h6ffff797;         'd997: data <= 32'h0b478793;
         'd998: data <= 32'h0007a403;         'd999: data <= 32'h00140413;
         'd1000: data <= 32'h0087a023;         'd1001: data <= 32'h04041c63;
         'd1002: data <= 32'h6ffff797;         'd1003: data <= 32'h0ac7a783;
         'd1004: data <= 32'h0007a783;         'd1005: data <= 32'h00078863;
         'd1006: data <= 32'h30047073;         'd1007: data <= 32'h00100073;
         'd1008: data <= 32'h0000006f;         'd1009: data <= 32'h6ffff717;
         'd1010: data <= 32'h09070713;         'd1011: data <= 32'h00072683;
         'd1012: data <= 32'h6ffff797;         'd1013: data <= 32'h08078793;
         'd1014: data <= 32'h0007a603;         'd1015: data <= 32'h00c72023;
         'd1016: data <= 32'h00d7a023;         'd1017: data <= 32'h6ffff717;
         'd1018: data <= 32'h04c70713;         'd1019: data <= 32'h00072783;
         'd1020: data <= 32'h00178793;         'd1021: data <= 32'h00f72023;
         'd1022: data <= 32'h819ff0ef;         'd1023: data <= 32'h6ffff797;
         'd1024: data <= 32'h02c7a783;         'd1025: data <= 32'h04f47e63;
         'd1026: data <= 32'h00000493;         'd1027: data <= 32'h6ffff797;
         'd1028: data <= 32'h04c7a783;         'd1029: data <= 32'h02c7a703;
         'd1030: data <= 32'h00271793;         'd1031: data <= 32'h00e787b3;
         'd1032: data <= 32'h00279713;         'd1033: data <= 32'h6ffff797;
         'd1034: data <= 32'h0e078793;         'd1035: data <= 32'h00e787b3;
         'd1036: data <= 32'h0007a703;         'd1037: data <= 32'h00100793;
         'd1038: data <= 32'h00e7f463;         'd1039: data <= 32'h00100493;
         'd1040: data <= 32'h6ffff797;         'd1041: data <= 32'hff87a783;
         'd1042: data <= 32'h16078e63;         'd1043: data <= 32'h6ffff797;
         'd1044: data <= 32'hfe87a783;         'd1045: data <= 32'h18078a63;
         'd1046: data <= 32'h00100493;         'd1047: data <= 32'h18c0006f;
         'd1048: data <= 32'h00000493;         'd1049: data <= 32'h0d00006f;
         'd1050: data <= 32'hfff00793;         'd1051: data <= 32'h6ffff717;
         'd1052: data <= 32'hfaf72e23;         'd1053: data <= 32'hf99ff06f;
         'd1054: data <= 32'h6ffff797;         'd1055: data <= 32'hfae7a823;
         'd1056: data <= 32'hf8dff06f;         'd1057: data <= 32'h00c7a683;
         'd1058: data <= 32'h00d72223;         'd1059: data <= 32'h0f40006f;
         'd1060: data <= 32'h0207a423;         'd1061: data <= 32'h00072683;
         'd1062: data <= 32'hfff68693;         'd1063: data <= 32'h00d72023;
         'd1064: data <= 32'h02c7a683;         'd1065: data <= 32'h00100713;
         'd1066: data <= 32'h00d71733;         'd1067: data <= 32'h6ffff617;
         'd1068: data <= 32'hf9460613;         'd1069: data <= 32'h00062503;
         'd1070: data <= 32'h00a76733;         'd1071: data <= 32'h00e62023;
         'd1072: data <= 32'h6ffff717;         'd1073: data <= 32'h04470713;
         'd1074: data <= 32'h00269613;         'd1075: data <= 32'h00d60633;
         'd1076: data <= 32'h00261693;         'd1077: data <= 32'h00d706b3;
         'd1078: data <= 32'h0046a683;         'd1079: data <= 32'h00d7a423;
         'd1080: data <= 32'h0086a603;         'd1081: data <= 32'h00c7a623;
         'd1082: data <= 32'h00b62223;         'd1083: data <= 32'h00b6a423;
         'd1084: data <= 32'h02c7a583;         'd1085: data <= 32'h00259693;
         'd1086: data <= 32'h00b68533;         'd1087: data <= 32'h00251613;
         'd1088: data <= 32'h00e60633;         'd1089: data <= 32'h00c7aa23;
         'd1090: data <= 32'h00062603;         'd1091: data <= 32'h00160613;
         'd1092: data <= 32'h00251593;         'd1093: data <= 32'h00b70733;
         'd1094: data <= 32'h00c72023;         'd1095: data <= 32'h02c7a703;
         'd1096: data <= 32'h6ffff797;         'd1097: data <= 32'hf387a783;
         'd1098: data <= 32'h02c7a783;         'd1099: data <= 32'h00f76463;
         'd1100: data <= 32'h00100493;         'd1101: data <= 32'h6ffff797;
         'd1102: data <= 32'hf207a783;         'd1103: data <= 32'h0007a783;
         'd1104: data <= 32'hf20784e3;         'd1105: data <= 32'h6ffff797;
         'd1106: data <= 32'hf107a783;         'd1107: data <= 32'h00c7a783;
         'd1108: data <= 32'h00c7a783;         'd1109: data <= 32'h0047a703;
         'd1110: data <= 32'hf2e460e3;         'd1111: data <= 32'h0147a703;
         'd1112: data <= 32'h0087a603;         'd1113: data <= 32'h00c7a683;
         'd1114: data <= 32'h00d62423;         'd1115: data <= 32'h0087a603;
         'd1116: data <= 32'h00c6a223;         'd1117: data <= 32'h00472683;
         'd1118: data <= 32'h00478593;         'd1119: data <= 32'hf0b684e3;
         'd1120: data <= 32'h0007aa23;         'd1121: data <= 32'h00072683;
         'd1122: data <= 32'hfff68693;         'd1123: data <= 32'h00d72023;
         'd1124: data <= 32'h0287a703;         'd1125: data <= 32'hf00706e3;
         'd1126: data <= 32'h01c7a603;         'd1127: data <= 32'h0207a683;
         'd1128: data <= 32'h00d62423;         'd1129: data <= 32'h01c7a603;
         'd1130: data <= 32'h00c6a223;         'd1131: data <= 32'h00472603;
         'd1132: data <= 32'h01878693;         'd1133: data <= 32'hecd61ee3;
         'd1134: data <= 32'h0207a683;         'd1135: data <= 32'h00d72223;
         'd1136: data <= 32'hed1ff06f;         'd1137: data <= 32'ha4cff0ef;
         'd1138: data <= 32'he85ff06f;         'd1139: data <= 32'h6ffff717;
         'd1140: data <= 32'he6c70713;         'd1141: data <= 32'h00072783;
         'd1142: data <= 32'h00178793;         'd1143: data <= 32'h00f72023;
         'd1144: data <= 32'ha30ff0ef;         'd1145: data <= 32'h00000493;
         'd1146: data <= 32'h00048513;         'd1147: data <= 32'h00c12083;
         'd1148: data <= 32'h00812403;         'd1149: data <= 32'h00412483;
         'd1150: data <= 32'h01010113;         'd1151: data <= 32'h00008067;
         'd1152: data <= 32'h6ffff797;         'd1153: data <= 32'he207a783;
         'd1154: data <= 32'h00079863;         'd1155: data <= 32'h30047073;
         'd1156: data <= 32'h00100073;         'd1157: data <= 32'h0000006f;
         'd1158: data <= 32'h30047073;         'd1159: data <= 32'h6ffff717;
         'd1160: data <= 32'hdf470713;         'd1161: data <= 32'h00072783;
         'd1162: data <= 32'h00178793;         'd1163: data <= 32'h00f72023;
         'd1164: data <= 32'h6ffff797;         'd1165: data <= 32'hdf078793;
         'd1166: data <= 32'h0007a703;         'd1167: data <= 32'hfff70713;
         'd1168: data <= 32'h00e7a023;         'd1169: data <= 32'h0007a783;
         'd1170: data <= 32'h1e079263;         'd1171: data <= 32'h6ffff797;
         'd1172: data <= 32'hdfc7a783;         'd1173: data <= 32'h02079263;
         'd1174: data <= 32'h00000513;         'd1175: data <= 32'h1d40006f;
         'd1176: data <= 32'h0207a683;         'd1177: data <= 32'h00d72223;
         'd1178: data <= 32'h05c0006f;         'd1179: data <= 32'h00c7a603;
         'd1180: data <= 32'h00c72223;         'd1181: data <= 32'h0840006f;
         'd1182: data <= 32'hff010113;         'd1183: data <= 32'h00112623;
         'd1184: data <= 32'h00812423;         'd1185: data <= 32'h00000793;
         'd1186: data <= 32'h6ffff717;         'd1187: data <= 32'he4072703;
         'd1188: data <= 32'h10070e63;         'd1189: data <= 32'h6ffff797;
         'd1190: data <= 32'he407a783;         'd1191: data <= 32'h00c7a783;
         'd1192: data <= 32'h0287a703;         'd1193: data <= 32'h01c7a603;
         'd1194: data <= 32'h0207a683;         'd1195: data <= 32'h00d62423;
         'd1196: data <= 32'h01c7a603;         'd1197: data <= 32'h00c6a223;
         'd1198: data <= 32'h00472603;         'd1199: data <= 32'h01878693;
         'd1200: data <= 32'hfad600e3;         'd1201: data <= 32'h0207a423;
         'd1202: data <= 32'h00072683;         'd1203: data <= 32'hfff68693;
         'd1204: data <= 32'h00d72023;         'd1205: data <= 32'h0147a703;
         'd1206: data <= 32'h0087a603;         'd1207: data <= 32'h00c7a683;
         'd1208: data <= 32'h00d62423;         'd1209: data <= 32'h0087a603;
         'd1210: data <= 32'h00c6a223;         'd1211: data <= 32'h00472603;
         'd1212: data <= 32'h00478693;         'd1213: data <= 32'hf6d60ce3;
         'd1214: data <= 32'h0007aa23;         'd1215: data <= 32'h00072603;
         'd1216: data <= 32'hfff60613;         'd1217: data <= 32'h00c72023;
         'd1218: data <= 32'h02c7a583;         'd1219: data <= 32'h00100713;
         'd1220: data <= 32'h00b71733;         'd1221: data <= 32'h6ffff617;
         'd1222: data <= 32'hd2c60613;         'd1223: data <= 32'h00062503;
         'd1224: data <= 32'h00a76733;         'd1225: data <= 32'h00e62023;
         'd1226: data <= 32'h6ffff617;         'd1227: data <= 32'hddc60613;
         'd1228: data <= 32'h00259713;         'd1229: data <= 32'h00b70733;
         'd1230: data <= 32'h00271713;         'd1231: data <= 32'h00e60733;
         'd1232: data <= 32'h00472703;         'd1233: data <= 32'h00e7a423;
         'd1234: data <= 32'h00872583;         'd1235: data <= 32'h00b7a623;
         'd1236: data <= 32'h00d5a223;         'd1237: data <= 32'h00d72423;
         'd1238: data <= 32'h02c7a583;         'd1239: data <= 32'h00259713;
         'd1240: data <= 32'h00b706b3;         'd1241: data <= 32'h00269693;
         'd1242: data <= 32'h00c686b3;         'd1243: data <= 32'h00d7aa23;
         'd1244: data <= 32'h0006a683;         'd1245: data <= 32'h00168693;
         'd1246: data <= 32'h00b70733;         'd1247: data <= 32'h00271713;
         'd1248: data <= 32'h00e60633;         'd1249: data <= 32'h00d62023;
         'd1250: data <= 32'h02c7a683;         'd1251: data <= 32'h6ffff717;
         'd1252: data <= 32'hccc72703;         'd1253: data <= 32'h02c72703;
         'd1254: data <= 32'heee6e8e3;         'd1255: data <= 32'h00100713;
         'd1256: data <= 32'h6ffff697;         'd1257: data <= 32'hc8e6aa23;
         'd1258: data <= 32'hee1ff06f;         'd1259: data <= 32'h00078463;
         'd1260: data <= 32'hc60ff0ef;         'd1261: data <= 32'h6ffff417;
         'd1262: data <= 32'hc8442403;         'd1263: data <= 32'h04041663;
         'd1264: data <= 32'h6ffff517;         'd1265: data <= 32'hc7452503;
         'd1266: data <= 32'h00050663;         'd1267: data <= 32'h00000073;
         'd1268: data <= 32'h00100513;         'd1269: data <= 32'h6ffff717;
         'd1270: data <= 32'hc3c70713;         'd1271: data <= 32'h00072783;
         'd1272: data <= 32'hfff78793;         'd1273: data <= 32'h00f72023;
         'd1274: data <= 32'h00079463;         'd1275: data <= 32'h30046073;
         'd1276: data <= 32'h00c12083;         'd1277: data <= 32'h00812403;
         'd1278: data <= 32'h01010113;         'd1279: data <= 32'h00008067;
         'd1280: data <= 32'hfff40413;         'd1281: data <= 32'h00040e63;
         'd1282: data <= 32'hb6dff0ef;         'd1283: data <= 32'hfe050ae3;
         'd1284: data <= 32'h00100793;         'd1285: data <= 32'h6ffff717;
         'd1286: data <= 32'hc2f72023;         'd1287: data <= 32'hfe5ff06f;
         'd1288: data <= 32'h6ffff797;         'd1289: data <= 32'hc007ac23;
         'd1290: data <= 32'hf99ff06f;         'd1291: data <= 32'h00000513;
         'd1292: data <= 32'h6ffff717;         'd1293: data <= 32'hbe070713;
         'd1294: data <= 32'h00072783;         'd1295: data <= 32'hfff78793;
         'd1296: data <= 32'h00f72023;         'd1297: data <= 32'h00079663;
         'd1298: data <= 32'h30046073;         'd1299: data <= 32'h00008067;
         'd1300: data <= 32'h00008067;         'd1301: data <= 32'h04050c63;
         'd1302: data <= 32'hff010113;         'd1303: data <= 32'h00112623;
         'd1304: data <= 32'h00812423;         'd1305: data <= 32'h00050413;
         'd1306: data <= 32'h6ffff797;         'd1307: data <= 32'hbb87a783;
         'd1308: data <= 32'h00078863;         'd1309: data <= 32'h30047073;
         'd1310: data <= 32'h00100073;         'd1311: data <= 32'h0000006f;
         'd1312: data <= 32'had1ff0ef;         'd1313: data <= 32'h00000593;
         'd1314: data <= 32'h00040513;         'd1315: data <= 32'hfecff0ef;
         'd1316: data <= 32'hd71ff0ef;         'd1317: data <= 32'h00051463;
         'd1318: data <= 32'h00000073;         'd1319: data <= 32'h00c12083;
         'd1320: data <= 32'h00812403;         'd1321: data <= 32'h01010113;
         'd1322: data <= 32'h00008067;         'd1323: data <= 32'h00000073;
         'd1324: data <= 32'h00008067;         'd1325: data <= 32'h6ffff797;
         'd1326: data <= 32'hb6c7a783;         'd1327: data <= 32'h00078a63;
         'd1328: data <= 32'h00100793;         'd1329: data <= 32'h6ffff717;
         'd1330: data <= 32'hb6f72823;         'd1331: data <= 32'h00008067;
         'd1332: data <= 32'hff010113;         'd1333: data <= 32'h00112623;
         'd1334: data <= 32'h6ffff797;         'd1335: data <= 32'hb407ae23;
         'd1336: data <= 32'h6ffff797;         'd1337: data <= 32'hb787a783;
         'd1338: data <= 32'h0307a703;         'd1339: data <= 32'h00072683;
         'd1340: data <= 32'ha5a5a7b7;         'd1341: data <= 32'h5a578793;
         'd1342: data <= 32'h00f69a63;         'd1343: data <= 32'h00472683;
         'd1344: data <= 32'ha5a5a7b7;         'd1345: data <= 32'h5a578793;
         'd1346: data <= 32'h04f68e63;         'd1347: data <= 32'h6ffff797;
         'd1348: data <= 32'hb4c78793;         'd1349: data <= 32'h0007a503;
         'd1350: data <= 32'h0007a583;         'd1351: data <= 32'h03458593;
         'd1352: data <= 32'hed1fe0ef;         'd1353: data <= 32'h6ffff517;
         'd1354: data <= 32'hb1c52503;         'd1355: data <= 32'h141010ef;
         'd1356: data <= 32'h01f00793;         'd1357: data <= 32'h40a78533;
         'd1358: data <= 32'h00251793;         'd1359: data <= 32'h00a787b3;
         'd1360: data <= 32'h00279793;         'd1361: data <= 32'h6ffff717;
         'd1362: data <= 32'hbc070713;         'd1363: data <= 32'h00f707b3;
         'd1364: data <= 32'h0007a783;         'd1365: data <= 32'h02079a63;
         'd1366: data <= 32'h30047073;         'd1367: data <= 32'h00100073;
         'd1368: data <= 32'h0000006f;         'd1369: data <= 32'h00872683;
         'd1370: data <= 32'ha5a5a7b7;         'd1371: data <= 32'h5a578793;
         'd1372: data <= 32'hf8f69ee3;         'd1373: data <= 32'h00c72703;
         'd1374: data <= 32'ha5a5a7b7;         'd1375: data <= 32'h5a578793;
         'd1376: data <= 32'hf8f716e3;         'd1377: data <= 32'hfa1ff06f;
         'd1378: data <= 32'h00251713;         'd1379: data <= 32'h00a70733;
         'd1380: data <= 32'h00271713;         'd1381: data <= 32'h6ffff797;
         'd1382: data <= 32'hb7078793;         'd1383: data <= 32'h00e787b3;
         'd1384: data <= 32'h0047a703;         'd1385: data <= 32'h00472703;
         'd1386: data <= 32'h00e7a223;         'd1387: data <= 32'h00878793;
         'd1388: data <= 32'h02f70c63;         'd1389: data <= 32'h00251793;
         'd1390: data <= 32'h00a787b3;         'd1391: data <= 32'h00279793;
         'd1392: data <= 32'h6ffff717;         'd1393: data <= 32'hb4470713;
         'd1394: data <= 32'h00f707b3;         'd1395: data <= 32'h0047a783;
         'd1396: data <= 32'h00c7a783;         'd1397: data <= 32'h6ffff717;
         'd1398: data <= 32'ha8f72223;         'd1399: data <= 32'h00c12083;
         'd1400: data <= 32'h01010113;         'd1401: data <= 32'h00008067;
         'd1402: data <= 32'h00472683;         'd1403: data <= 32'h00251793;
         'd1404: data <= 32'h00a787b3;         'd1405: data <= 32'h00279793;
         'd1406: data <= 32'h6ffff717;         'd1407: data <= 32'hb0c70713;
         'd1408: data <= 32'h00f707b3;         'd1409: data <= 32'h00d7a223;
         'd1410: data <= 32'hfadff06f;         'd1411: data <= 32'h04050063;
         'd1412: data <= 32'hff010113;         'd1413: data <= 32'h00112623;
         'd1414: data <= 32'h00812423;         'd1415: data <= 32'h00058413;
         'd1416: data <= 32'h6ffff597;         'd1417: data <= 32'ha385a583;
         'd1418: data <= 32'h01858593;         'd1419: data <= 32'h505000ef;
         'd1420: data <= 32'h00100593;         'd1421: data <= 32'h00040513;
         'd1422: data <= 32'he40ff0ef;         'd1423: data <= 32'h00c12083;
         'd1424: data <= 32'h00812403;         'd1425: data <= 32'h01010113;
         'd1426: data <= 32'h00008067;         'd1427: data <= 32'h30047073;
         'd1428: data <= 32'h00100073;         'd1429: data <= 32'h0000006f;
         'd1430: data <= 32'h00050793;         'd1431: data <= 32'h06050c63;
         'd1432: data <= 32'hff010113;         'd1433: data <= 32'h00112623;
         'd1434: data <= 32'h00058513;         'd1435: data <= 32'h00060593;
         'd1436: data <= 32'h0047a683;         'd1437: data <= 32'h6ffff717;
         'd1438: data <= 32'h9e470713;         'd1439: data <= 32'h00072603;
         'd1440: data <= 32'h00d62e23;         'd1441: data <= 32'h00072603;
         'd1442: data <= 32'h0086a803;         'd1443: data <= 32'h03062023;
         'd1444: data <= 32'h00072603;         'd1445: data <= 32'h01860613;
         'd1446: data <= 32'h00c82223;         'd1447: data <= 32'h00072603;
         'd1448: data <= 32'h01860613;         'd1449: data <= 32'h00c6a423;
         'd1450: data <= 32'h00072703;         'd1451: data <= 32'h02f72423;
         'd1452: data <= 32'h0007a703;         'd1453: data <= 32'h00170713;
         'd1454: data <= 32'h00e7a023;         'd1455: data <= 32'h00058463;
         'd1456: data <= 32'hfff00513;         'd1457: data <= 32'hdb4ff0ef;
         'd1458: data <= 32'h00c12083;         'd1459: data <= 32'h01010113;
         'd1460: data <= 32'h00008067;         'd1461: data <= 32'h30047073;
         'd1462: data <= 32'h00100073;         'd1463: data <= 32'h0000006f;
         'd1464: data <= 32'h00c52783;         'd1465: data <= 32'h00c7a783;
         'd1466: data <= 32'h12078063;         'd1467: data <= 32'h0287a703;
         'd1468: data <= 32'h01c7a603;         'd1469: data <= 32'h0207a683;
         'd1470: data <= 32'h00d62423;         'd1471: data <= 32'h01c7a603;
         'd1472: data <= 32'h00c6a223;         'd1473: data <= 32'h00472683;
         'd1474: data <= 32'h01878613;         'd1475: data <= 32'h10c68463;
         'd1476: data <= 32'h0207a423;         'd1477: data <= 32'h00072683;
         'd1478: data <= 32'hfff68693;         'd1479: data <= 32'h00d72023;
         'd1480: data <= 32'h6ffff717;         'd1481: data <= 32'h90072703;
         'd1482: data <= 32'h10071263;         'd1483: data <= 32'h0147a703;
         'd1484: data <= 32'h0087a603;         'd1485: data <= 32'h00c7a683;
         'd1486: data <= 32'h00d62423;         'd1487: data <= 32'h0087a603;
         'd1488: data <= 32'h00c6a223;         'd1489: data <= 32'h00472603;
         'd1490: data <= 32'h00478693;         'd1491: data <= 32'h0cd60a63;
         'd1492: data <= 32'h0007aa23;         'd1493: data <= 32'h00072603;
         'd1494: data <= 32'hfff60613;         'd1495: data <= 32'h00c72023;
         'd1496: data <= 32'h02c7a583;         'd1497: data <= 32'h00100713;
         'd1498: data <= 32'h00b71733;         'd1499: data <= 32'h6ffff617;
         'd1500: data <= 32'h8d460613;         'd1501: data <= 32'h00062503;
         'd1502: data <= 32'h00a76733;         'd1503: data <= 32'h00e62023;
         'd1504: data <= 32'h6ffff617;         'd1505: data <= 32'h98460613;
         'd1506: data <= 32'h00259713;         'd1507: data <= 32'h00b70733;
         'd1508: data <= 32'h00271713;         'd1509: data <= 32'h00e60733;
         'd1510: data <= 32'h00472703;         'd1511: data <= 32'h00e7a423;
         'd1512: data <= 32'h00872583;         'd1513: data <= 32'h00b7a623;
         'd1514: data <= 32'h00d5a223;         'd1515: data <= 32'h00d72423;
         'd1516: data <= 32'h02c7a583;         'd1517: data <= 32'h00259713;
         'd1518: data <= 32'h00b706b3;         'd1519: data <= 32'h00269693;
         'd1520: data <= 32'h00c686b3;         'd1521: data <= 32'h00d7aa23;
         'd1522: data <= 32'h0006a683;         'd1523: data <= 32'h00168693;
         'd1524: data <= 32'h00b70733;         'd1525: data <= 32'h00271713;
         'd1526: data <= 32'h00e60633;         'd1527: data <= 32'h00d62023;
         'd1528: data <= 32'h02c7a703;         'd1529: data <= 32'h6ffff797;
         'd1530: data <= 32'h8747a783;         'd1531: data <= 32'h02c7a783;
         'd1532: data <= 32'h06e7f863;         'd1533: data <= 32'h00100793;
         'd1534: data <= 32'h6ffff717;         'd1535: data <= 32'h82f72e23;
         'd1536: data <= 32'h00100513;         'd1537: data <= 32'h00008067;
         'd1538: data <= 32'h30047073;         'd1539: data <= 32'h00100073;
         'd1540: data <= 32'h0000006f;         'd1541: data <= 32'h0207a683;
         'd1542: data <= 32'h00d72223;         'd1543: data <= 32'hef5ff06f;
         'd1544: data <= 32'h00c7a603;         'd1545: data <= 32'h00c72223;
         'd1546: data <= 32'hf29ff06f;         'd1547: data <= 32'h6ffff717;
         'd1548: data <= 32'h89c70713;         'd1549: data <= 32'h00472683;
         'd1550: data <= 32'h00d7ae23;         'd1551: data <= 32'h0086a583;
         'd1552: data <= 32'h02b7a023;         'd1553: data <= 32'h00c5a223;
         'd1554: data <= 32'h00c6a423;         'd1555: data <= 32'h02e7a423;
         'd1556: data <= 32'h00072683;         'd1557: data <= 32'h00168693;
         'd1558: data <= 32'h00d72023;         'd1559: data <= 32'hf85ff06f;
         'd1560: data <= 32'h00000513;         'd1561: data <= 32'h00008067;
         'd1562: data <= 32'h6fffe797;         'd1563: data <= 32'h7c87a783;
         'd1564: data <= 32'h00f52023;         'd1565: data <= 32'h6fffe797;
         'd1566: data <= 32'h7d07a783;         'd1567: data <= 32'h00f52223;
         'd1568: data <= 32'h00008067;         'd1569: data <= 32'h06050863;
         'd1570: data <= 32'h06058c63;         'd1571: data <= 32'h30047073;
         'd1572: data <= 32'h6fffe717;         'd1573: data <= 32'h78070713;
         'd1574: data <= 32'h00072783;         'd1575: data <= 32'h00178793;
         'd1576: data <= 32'h00f72023;         'd1577: data <= 32'h6fffe717;
         'd1578: data <= 32'h7a072703;         'd1579: data <= 32'h00452783;
         'd1580: data <= 32'h40f70633;         'd1581: data <= 32'h6fffe697;
         'd1582: data <= 32'h7a46a683;         'd1583: data <= 32'h0606c683;
         'd1584: data <= 32'h04068663;         'd1585: data <= 32'h6fffe797;
         'd1586: data <= 32'h7947a783;         'd1587: data <= 32'h06078023;
         'd1588: data <= 32'h00100513;         'd1589: data <= 32'h6fffe717;
         'd1590: data <= 32'h73c70713;         'd1591: data <= 32'h00072783;
         'd1592: data <= 32'hfff78793;         'd1593: data <= 32'h00f72023;
         'd1594: data <= 32'h0a079663;         'd1595: data <= 32'h30046073;
         'd1596: data <= 32'h00008067;         'd1597: data <= 32'h30047073;
         'd1598: data <= 32'h00100073;         'd1599: data <= 32'h0000006f;
         'd1600: data <= 32'h30047073;         'd1601: data <= 32'h00100073;
         'd1602: data <= 32'h0000006f;         'd1603: data <= 32'h0005a683;
         'd1604: data <= 32'hfff00813;         'd1605: data <= 32'h03068a63;
         'd1606: data <= 32'h00052883;         'd1607: data <= 32'h6fffe817;
         'd1608: data <= 32'h71482803;         'd1609: data <= 32'h01088a63;
         'd1610: data <= 32'h00f76863;         'd1611: data <= 32'h0005a023;
         'd1612: data <= 32'h00100513;         'd1613: data <= 32'hfa1ff06f;
         'd1614: data <= 32'h00d66c63;         'd1615: data <= 32'h0005a023;
         'd1616: data <= 32'h00100513;         'd1617: data <= 32'hf91ff06f;
         'd1618: data <= 32'h00000513;         'd1619: data <= 32'hf89ff06f;
         'd1620: data <= 32'hff010113;         'd1621: data <= 32'h00112623;
         'd1622: data <= 32'h40e787b3;         'd1623: data <= 32'h00d787b3;
         'd1624: data <= 32'h00f5a023;         'd1625: data <= 32'hf05ff0ef;
         'd1626: data <= 32'h00000513;         'd1627: data <= 32'h6fffe717;
         'd1628: data <= 32'h6a470713;         'd1629: data <= 32'h00072783;
         'd1630: data <= 32'hfff78793;         'd1631: data <= 32'h00f72023;
         'd1632: data <= 32'h00079463;         'd1633: data <= 32'h30046073;
         'd1634: data <= 32'h00c12083;         'd1635: data <= 32'h01010113;
         'd1636: data <= 32'h00008067;         'd1637: data <= 32'h00008067;
         'd1638: data <= 32'h00100793;         'd1639: data <= 32'h6fffe717;
         'd1640: data <= 32'h68f72c23;         'd1641: data <= 32'h00008067;
         'd1642: data <= 32'h6fffe797;         'd1643: data <= 32'h6947a783;
         'd1644: data <= 32'h02078063;         'd1645: data <= 32'h6fffe797;
         'd1646: data <= 32'h66c7a783;         'd1647: data <= 32'h00078663;
         'd1648: data <= 32'h00000513;         'd1649: data <= 32'h00008067;
         'd1650: data <= 32'h00200513;         'd1651: data <= 32'h00008067;
         'd1652: data <= 32'h00100513;         'd1653: data <= 32'h00008067;
         'd1654: data <= 32'h6fffe717;         'd1655: data <= 32'h69472703;
         'd1656: data <= 32'h00072783;         'd1657: data <= 32'h00079e63;
         'd1658: data <= 32'h00100793;         'd1659: data <= 32'h00f52023;
         'd1660: data <= 32'h00079c63;         'd1661: data <= 32'h00c72783;
         'd1662: data <= 32'h0007a503;         'd1663: data <= 32'h00008067;
         'd1664: data <= 32'h00000793;         'd1665: data <= 32'hfe9ff06f;
         'd1666: data <= 32'h00000513;         'd1667: data <= 32'h00008067;
         'd1668: data <= 32'hff010113;         'd1669: data <= 32'h00112623;
         'd1670: data <= 32'h00b52223;         'd1671: data <= 32'h00a52823;
         'd1672: data <= 32'h02b66c63;         'd1673: data <= 32'h40d60633;
         'd1674: data <= 32'h01852783;         'd1675: data <= 32'h00f66a63;
         'd1676: data <= 32'h00100513;         'd1677: data <= 32'h00c12083;
         'd1678: data <= 32'h01010113;         'd1679: data <= 32'h00008067;
         'd1680: data <= 32'h00450593;         'd1681: data <= 32'h6fffe517;
         'd1682: data <= 32'h62452503;         'd1683: data <= 32'h0e5000ef;
         'd1684: data <= 32'h00000513;         'd1685: data <= 32'hfe1ff06f;
         'd1686: data <= 32'h00d67463;         'd1687: data <= 32'h00d5fe63;
         'd1688: data <= 32'h00450593;         'd1689: data <= 32'h6fffe517;
         'd1690: data <= 32'h60852503;         'd1691: data <= 32'h0c5000ef;
         'd1692: data <= 32'h00000513;         'd1693: data <= 32'hfc1ff06f;
         'd1694: data <= 32'h00100513;         'd1695: data <= 32'hfb9ff06f;
         'd1696: data <= 32'hff010113;         'd1697: data <= 32'h00112623;
         'd1698: data <= 32'h00812423;         'd1699: data <= 32'h00912223;
         'd1700: data <= 32'h01212023;         'd1701: data <= 32'h00050413;
         'd1702: data <= 32'h00058493;         'd1703: data <= 32'h00060913;
         'd1704: data <= 32'h0180006f;         'd1705: data <= 32'h01842783;
         'd1706: data <= 32'h00f484b3;         'd1707: data <= 32'h02042783;
         'd1708: data <= 32'h00040513;         'd1709: data <= 32'h000780e7;
         'd1710: data <= 32'h01842583;         'd1711: data <= 32'h00048693;
         'd1712: data <= 32'h00090613;         'd1713: data <= 32'h009585b3;
         'd1714: data <= 32'h00040513;         'd1715: data <= 32'hf45ff0ef;
         'd1716: data <= 32'hfc051ae3;         'd1717: data <= 32'h00c12083;
         'd1718: data <= 32'h00812403;         'd1719: data <= 32'h00412483;
         'd1720: data <= 32'h00012903;         'd1721: data <= 32'h01010113;
         'd1722: data <= 32'h00008067;         'd1723: data <= 32'hff010113;
         'd1724: data <= 32'h00112623;         'd1725: data <= 32'h00812423;
         'd1726: data <= 32'h00912223;         'd1727: data <= 32'h01212023;
         'd1728: data <= 32'h00050493;         'd1729: data <= 32'h00058913;
         'd1730: data <= 32'h6fffe797;         'd1731: data <= 32'h5647a783;
         'd1732: data <= 32'h00c7a783;         'd1733: data <= 32'h00c7a403;
         'd1734: data <= 32'h00440513;         'd1735: data <= 32'h065000ef;
         'd1736: data <= 32'h02444783;         'd1737: data <= 32'h0047f713;
         'd1738: data <= 32'h02071863;         'd1739: data <= 32'hffe7f793;
         'd1740: data <= 32'h02f40223;         'd1741: data <= 32'h02042783;
         'd1742: data <= 32'h00040513;         'd1743: data <= 32'h000780e7;
         'd1744: data <= 32'h00c12083;         'd1745: data <= 32'h00812403;
         'd1746: data <= 32'h00412483;         'd1747: data <= 32'h00012903;
         'd1748: data <= 32'h01010113;         'd1749: data <= 32'h00008067;
         'd1750: data <= 32'h00090613;         'd1751: data <= 32'h00048593;
         'd1752: data <= 32'h00040513;         'd1753: data <= 32'hf1dff0ef;
         'd1754: data <= 32'hfcdff06f;         'd1755: data <= 32'h6fffe797;
         'd1756: data <= 32'h5007a783;         'd1757: data <= 32'h0007a703;
         'd1758: data <= 32'h04070863;         'd1759: data <= 32'hff010113;
         'd1760: data <= 32'h00112623;         'd1761: data <= 32'h00c7a783;
         'd1762: data <= 32'hfff00593;         'd1763: data <= 32'h0007a503;
         'd1764: data <= 32'hf5dff0ef;         'd1765: data <= 32'h6fffe797;
         'd1766: data <= 32'h4d87a783;         'd1767: data <= 32'h0007a703;
         'd1768: data <= 32'hfe0712e3;         'd1769: data <= 32'h6fffe717;
         'd1770: data <= 32'h4c470713;         'd1771: data <= 32'h00072683;
         'd1772: data <= 32'h6fffe617;         'd1773: data <= 32'h4ad62e23;
         'd1774: data <= 32'h00f72023;         'd1775: data <= 32'h00c12083;
         'd1776: data <= 32'h01010113;         'd1777: data <= 32'h00008067;
         'd1778: data <= 32'h6fffe717;         'd1779: data <= 32'h4a070713;
         'd1780: data <= 32'h00072683;         'd1781: data <= 32'h6fffe617;
         'd1782: data <= 32'h48d62c23;         'd1783: data <= 32'h00f72023;
         'd1784: data <= 32'h00008067;         'd1785: data <= 32'hff010113;
         'd1786: data <= 32'h00112623;         'd1787: data <= 32'h00812423;
         'd1788: data <= 32'h00912223;         'd1789: data <= 32'h00050493;
         'd1790: data <= 32'hb70ff0ef;         'd1791: data <= 32'h00050413;
         'd1792: data <= 32'h6fffe797;         'd1793: data <= 32'h45c7a783;
         'd1794: data <= 32'h02f56463;         'd1795: data <= 32'h0004a023;
         'd1796: data <= 32'h6fffe797;         'd1797: data <= 32'h4487a623;
         'd1798: data <= 32'h00040513;         'd1799: data <= 32'h00c12083;
         'd1800: data <= 32'h00812403;         'd1801: data <= 32'h00412483;
         'd1802: data <= 32'h01010113;         'd1803: data <= 32'h00008067;
         'd1804: data <= 32'hf3dff0ef;         'd1805: data <= 32'h00100793;
         'd1806: data <= 32'h00f4a023;         'd1807: data <= 32'hfd5ff06f;
         'd1808: data <= 32'hfe010113;         'd1809: data <= 32'h00112e23;
         'd1810: data <= 32'h00812c23;         'd1811: data <= 32'h00912a23;
         'd1812: data <= 32'h01212823;         'd1813: data <= 32'h00050913;
         'd1814: data <= 32'h00058413;         'd1815: data <= 32'haf4ff0ef;
         'd1816: data <= 32'h00c10513;         'd1817: data <= 32'hf81ff0ef;
         'd1818: data <= 32'h00c12783;         'd1819: data <= 32'h06079463;
         'd1820: data <= 32'h00050493;         'd1821: data <= 32'h04041063;
         'd1822: data <= 32'h03257463;         'd1823: data <= 32'h00040613;
         'd1824: data <= 32'h409905b3;         'd1825: data <= 32'h6fffe517;
         'd1826: data <= 32'h3e052503;         'd1827: data <= 32'h6c5000ef;
         'd1828: data <= 32'hd70ff0ef;         'd1829: data <= 32'h04051263;
         'd1830: data <= 32'h00000073;         'd1831: data <= 32'h03c0006f;
         'd1832: data <= 32'hd60ff0ef;         'd1833: data <= 32'h00048593;
         'd1834: data <= 32'h00090513;         'd1835: data <= 32'he41ff0ef;
         'd1836: data <= 32'h0280006f;         'd1837: data <= 32'h6fffe717;
         'd1838: data <= 32'h3b472703;         'd1839: data <= 32'h00072703;
         'd1840: data <= 32'h00071663;         'd1841: data <= 32'h00100413;
         'd1842: data <= 32'hfb5ff06f;         'd1843: data <= 32'h00078413;
         'd1844: data <= 32'hfadff06f;         'd1845: data <= 32'hd2cff0ef;
         'd1846: data <= 32'h01c12083;         'd1847: data <= 32'h01812403;
         'd1848: data <= 32'h01412483;         'd1849: data <= 32'h01012903;
         'd1850: data <= 32'h02010113;         'd1851: data <= 32'h00008067;
         'd1852: data <= 32'hfd010113;         'd1853: data <= 32'h02112623;
         'd1854: data <= 32'h02812423;         'd1855: data <= 32'h02912223;
         'd1856: data <= 32'h00c0006f;         'd1857: data <= 32'h01012783;
         'd1858: data <= 32'h0207dc63;         'd1859: data <= 32'h00000613;
         'd1860: data <= 32'h01010593;         'd1861: data <= 32'h6fffe517;
         'd1862: data <= 32'h35052503;         'd1863: data <= 32'h37d000ef;
         'd1864: data <= 32'h14050063;         'd1865: data <= 32'h01012783;
         'd1866: data <= 32'hfc07dee3;         'd1867: data <= 32'h01c12583;
         'd1868: data <= 32'h01812503;         'd1869: data <= 32'h01412783;
         'd1870: data <= 32'h000780e7;         'd1871: data <= 32'hfc9ff06f;
         'd1872: data <= 32'h01812403;         'd1873: data <= 32'h01442783;
         'd1874: data <= 32'h00078663;         'd1875: data <= 32'h00440513;
         'd1876: data <= 32'h630000ef;         'd1877: data <= 32'h00c10513;
         'd1878: data <= 32'he8dff0ef;         'd1879: data <= 32'h00050493;
         'd1880: data <= 32'h01012783;         'd1881: data <= 32'h00900713;
         'd1882: data <= 32'hfaf762e3;         'd1883: data <= 32'h00279793;
         'd1884: data <= 32'h00002717;         'd1885: data <= 32'h8b070713;
         'd1886: data <= 32'h00e787b3;         'd1887: data <= 32'h0007a783;
         'd1888: data <= 32'h00e787b3;         'd1889: data <= 32'h00078067;
         'd1890: data <= 32'h02444783;         'd1891: data <= 32'h0017e793;
         'd1892: data <= 32'h02f40223;         'd1893: data <= 32'h01412683;
         'd1894: data <= 32'h01842583;         'd1895: data <= 32'h00050613;
         'd1896: data <= 32'h00b685b3;         'd1897: data <= 32'h00040513;
         'd1898: data <= 32'hc69ff0ef;         'd1899: data <= 32'hf60500e3;
         'd1900: data <= 32'h02444783;         'd1901: data <= 32'h0047f713;
         'd1902: data <= 32'h00071e63;         'd1903: data <= 32'hffe7f793;
         'd1904: data <= 32'h02f40223;         'd1905: data <= 32'h02042783;
         'd1906: data <= 32'h00040513;         'd1907: data <= 32'h000780e7;
         'd1908: data <= 32'hf3dff06f;         'd1909: data <= 32'h01842783;
         'd1910: data <= 32'h00048613;         'd1911: data <= 32'h01412583;
         'd1912: data <= 32'h00f585b3;         'd1913: data <= 32'h00040513;
         'd1914: data <= 32'hc99ff0ef;         'd1915: data <= 32'hfd9ff06f;
         'd1916: data <= 32'h02444783;         'd1917: data <= 32'hffe7f793;
         'd1918: data <= 32'h02f40223;         'd1919: data <= 32'hf11ff06f;
         'd1920: data <= 32'h02444783;         'd1921: data <= 32'h0017e793;
         'd1922: data <= 32'h02f40223;         'd1923: data <= 32'h01412583;
         'd1924: data <= 32'h00b42c23;         'd1925: data <= 32'h00058e63;
         'd1926: data <= 32'h00050693;         'd1927: data <= 32'h00050613;
         'd1928: data <= 32'h00a585b3;         'd1929: data <= 32'h00040513;
         'd1930: data <= 32'hbe9ff0ef;         'd1931: data <= 32'hee1ff06f;
         'd1932: data <= 32'h30047073;         'd1933: data <= 32'h00100073;
         'd1934: data <= 32'h0000006f;         'd1935: data <= 32'h02444783;
         'd1936: data <= 32'h0027f713;         'd1937: data <= 32'h00070863;
         'd1938: data <= 32'hffe7f793;         'd1939: data <= 32'h02f40223;
         'd1940: data <= 32'hebdff06f;         'd1941: data <= 32'h00040513;
         'd1942: data <= 32'h400000ef;         'd1943: data <= 32'heb1ff06f;
         'd1944: data <= 32'h02c12083;         'd1945: data <= 32'h02812403;
         'd1946: data <= 32'h02412483;         'd1947: data <= 32'h03010113;
         'd1948: data <= 32'h00008067;         'd1949: data <= 32'hfe010113;
         'd1950: data <= 32'h00112e23;         'd1951: data <= 32'h00c10513;
         'd1952: data <= 32'hb59ff0ef;         'd1953: data <= 32'h00c12583;
         'd1954: data <= 32'hdb9ff0ef;         'd1955: data <= 32'he65ff0ef;
         'd1956: data <= 32'hfedff06f;         'd1957: data <= 32'h30047073;
         'd1958: data <= 32'h6fffe717;         'd1959: data <= 32'h17870713;
         'd1960: data <= 32'h00072783;         'd1961: data <= 32'h00178793;
         'd1962: data <= 32'h00f72023;         'd1963: data <= 32'h6fffe797;
         'd1964: data <= 32'h1b87a783;         'd1965: data <= 32'h02078263;
         'd1966: data <= 32'h6fffe717;         'd1967: data <= 32'h15870713;
         'd1968: data <= 32'h00072783;         'd1969: data <= 32'hfff78793;
         'd1970: data <= 32'h00f72023;         'd1971: data <= 32'h08079663;
         'd1972: data <= 32'h30046073;         'd1973: data <= 32'h00008067;
         'd1974: data <= 32'hff010113;         'd1975: data <= 32'h00112623;
         'd1976: data <= 32'h96418513;         'd1977: data <= 32'h424000ef;
         'd1978: data <= 32'h95018513;         'd1979: data <= 32'h41c000ef;
         'd1980: data <= 32'h96418793;         'd1981: data <= 32'h6fffe717;
         'd1982: data <= 32'h16f72c23;         'd1983: data <= 32'h95018793;
         'd1984: data <= 32'h6fffe717;         'd1985: data <= 32'h16f72423;
         'd1986: data <= 32'h00000613;         'd1987: data <= 32'h01000593;
         'd1988: data <= 32'h00400513;         'd1989: data <= 32'h04d000ef;
         'd1990: data <= 32'h6fffe797;         'd1991: data <= 32'h14a7a623;
         'd1992: data <= 32'h00050863;         'd1993: data <= 32'h00001597;
         'd1994: data <= 32'h72458593;         'd1995: data <= 32'h391000ef;
         'd1996: data <= 32'h6fffe717;         'd1997: data <= 32'h0e070713;
         'd1998: data <= 32'h00072783;         'd1999: data <= 32'hfff78793;
         'd2000: data <= 32'h00f72023;         'd2001: data <= 32'h00079463;
         'd2002: data <= 32'h30046073;         'd2003: data <= 32'h00c12083;
         'd2004: data <= 32'h01010113;         'd2005: data <= 32'h00008067;
         'd2006: data <= 32'h00008067;         'd2007: data <= 32'hff010113;
         'd2008: data <= 32'h00112623;         'd2009: data <= 32'hf31ff0ef;
         'd2010: data <= 32'h6fffe797;         'd2011: data <= 32'h0fc7a783;
         'd2012: data <= 32'h02078863;         'd2013: data <= 32'h6fffe797;
         'd2014: data <= 32'h0ec78793;         'd2015: data <= 32'h00400713;
         'd2016: data <= 32'h00000693;         'd2017: data <= 32'h08000613;
         'd2018: data <= 32'h00001597;         'd2019: data <= 32'h6c858593;
         'd2020: data <= 32'h00000517;         'd2021: data <= 32'hee450513;
         'd2022: data <= 32'he3dfe0ef;         'd2023: data <= 32'h00051863;
         'd2024: data <= 32'h30047073;         'd2025: data <= 32'h00100073;
         'd2026: data <= 32'h0000006f;         'd2027: data <= 32'h00c12083;
         'd2028: data <= 32'h01010113;         'd2029: data <= 32'h00008067;
         'd2030: data <= 32'h6fffe717;         'd2031: data <= 32'h1d870713;
         'd2032: data <= 32'h00f77793;         'd2033: data <= 32'h06078863;
         'd2034: data <= 32'h6fffe697;         'd2035: data <= 32'h1d768693;
         'd2036: data <= 32'hff06f693;         'd2037: data <= 32'h000027b7;
         'd2038: data <= 32'hc0078793;         'd2039: data <= 32'h40d787b3;
         'd2040: data <= 32'h00e787b3;         'd2041: data <= 32'h00068713;
         'd2042: data <= 32'h6fffe697;         'd2043: data <= 32'h09c68693;
         'd2044: data <= 32'h00e6a023;         'd2045: data <= 32'h0006a223;
         'd2046: data <= 32'h00f707b3;         'd2047: data <= 32'hff078793;
         'd2048: data <= 32'hff07f793;         'd2049: data <= 32'h6fffe697;
         'd2050: data <= 32'h06f6ae23;         'd2051: data <= 32'h0007a223;
         'd2052: data <= 32'h0007a023;         'd2053: data <= 32'h40e786b3;
         'd2054: data <= 32'h00d72223;         'd2055: data <= 32'h00f72023;
         'd2056: data <= 32'h6fffe797;         'd2057: data <= 32'h04d7ac23;
         'd2058: data <= 32'h6fffe797;         'd2059: data <= 32'h04d7aa23;
         'd2060: data <= 32'h00008067;         'd2061: data <= 32'h000027b7;
         'd2062: data <= 32'hc0078793;         'd2063: data <= 32'hfadff06f;
         'd2064: data <= 32'h6fffe797;         'd2065: data <= 32'h04478793;
         'd2066: data <= 32'h00078713;         'd2067: data <= 32'h0007a783;
         'd2068: data <= 32'hfea7ece3;         'd2069: data <= 32'h00472683;
         'd2070: data <= 32'h00d70633;         'd2071: data <= 32'h02a60063;
         'd2072: data <= 32'h00452683;         'd2073: data <= 32'h00d50633;
         'd2074: data <= 32'h02c78463;         'd2075: data <= 32'h00f52023;
         'd2076: data <= 32'h00e50463;         'd2077: data <= 32'h00a72023;
         'd2078: data <= 32'h00008067;         'd2079: data <= 32'h00452603;
         'd2080: data <= 32'h00c686b3;         'd2081: data <= 32'h00d72223;
         'd2082: data <= 32'h00070513;         'd2083: data <= 32'hfd5ff06f;
         'd2084: data <= 32'h6fffe617;         'd2085: data <= 32'hff062603;
         'd2086: data <= 32'h02c78063;         'd2087: data <= 32'h0047a783;
         'd2088: data <= 32'h00f686b3;         'd2089: data <= 32'h00d52223;
         'd2090: data <= 32'h00072783;         'd2091: data <= 32'h0007a783;
         'd2092: data <= 32'h00f52023;         'd2093: data <= 32'hfbdff06f;
         'd2094: data <= 32'h00c52023;         'd2095: data <= 32'hfb5ff06f;
         'd2096: data <= 32'hff010113;         'd2097: data <= 32'h00112623;
         'd2098: data <= 32'h00812423;         'd2099: data <= 32'h00912223;
         'd2100: data <= 32'h01212023;         'd2101: data <= 32'h00050493;
         'd2102: data <= 32'he79fe0ef;         'd2103: data <= 32'h6fffe797;
         'd2104: data <= 32'hfa47a783;         'd2105: data <= 32'h02078863;
         'd2106: data <= 32'h02048c63;         'd2107: data <= 32'h00f4f793;
         'd2108: data <= 32'h02000713;         'd2109: data <= 32'h40f70733;
         'd2110: data <= 32'hfdf78793;         'd2111: data <= 32'h0297e063;
         'd2112: data <= 32'h00e484b3;         'd2113: data <= 32'h0004de63;
         'd2114: data <= 32'h8f8ff0ef;         'd2115: data <= 32'h00000913;
         'd2116: data <= 32'h0380006f;         'd2117: data <= 32'hea5ff0ef;
         'd2118: data <= 32'hfd1ff06f;         'd2119: data <= 32'h00000493;
         'd2120: data <= 32'h02048063;         'd2121: data <= 32'h6fffe797;
         'd2122: data <= 32'hf587a783;         'd2123: data <= 32'h0297ea63;
         'd2124: data <= 32'h6fffe717;         'd2125: data <= 32'hf5470713;
         'd2126: data <= 32'h00072403;         'd2127: data <= 32'h0380006f;
         'd2128: data <= 32'h8c0ff0ef;         'd2129: data <= 32'h00000913;
         'd2130: data <= 32'ha84fe0ef;         'd2131: data <= 32'h00f97793;
         'd2132: data <= 32'h0e078663;         'd2133: data <= 32'h30047073;
         'd2134: data <= 32'h00100073;         'd2135: data <= 32'h0000006f;
         'd2136: data <= 32'h8a0ff0ef;         'd2137: data <= 32'h00000913;
         'd2138: data <= 32'hfe1ff06f;         'd2139: data <= 32'h00040713;
         'd2140: data <= 32'h00078413;         'd2141: data <= 32'h00442783;
         'd2142: data <= 32'h0097f663;         'd2143: data <= 32'h00042783;
         'd2144: data <= 32'hfe0796e3;         'd2145: data <= 32'h6fffe797;
         'd2146: data <= 32'hefc7a783;         'd2147: data <= 32'h02878e63;
         'd2148: data <= 32'h00072903;         'd2149: data <= 32'h01090913;
         'd2150: data <= 32'h00042783;         'd2151: data <= 32'h00f72023;
         'd2152: data <= 32'h00442783;         'd2153: data <= 32'h409787b3;
         'd2154: data <= 32'h02000713;         'd2155: data <= 32'h02f77a63;
         'd2156: data <= 32'h00940533;         'd2157: data <= 32'h00f57713;
         'd2158: data <= 32'h00070e63;         'd2159: data <= 32'h30047073;
         'd2160: data <= 32'h00100073;         'd2161: data <= 32'h0000006f;
         'd2162: data <= 32'h838ff0ef;         'd2163: data <= 32'h00000913;
         'd2164: data <= 32'hf79ff06f;         'd2165: data <= 32'h00f52223;
         'd2166: data <= 32'h00942223;         'd2167: data <= 32'he65ff0ef;
         'd2168: data <= 32'h00442703;         'd2169: data <= 32'h6fffe697;
         'd2170: data <= 32'he9868693;         'd2171: data <= 32'h0006a783;
         'd2172: data <= 32'h40e787b3;         'd2173: data <= 32'h00f6a023;
         'd2174: data <= 32'h6fffe697;         'd2175: data <= 32'he806a683;
         'd2176: data <= 32'h00d7f663;         'd2177: data <= 32'h6fffe697;
         'd2178: data <= 32'he6f6aa23;         'd2179: data <= 32'h800007b7;
         'd2180: data <= 32'h00f76733;         'd2181: data <= 32'h00e42223;
         'd2182: data <= 32'h00042023;         'd2183: data <= 32'h6fffe717;
         'd2184: data <= 32'he5870713;         'd2185: data <= 32'h00072783;
         'd2186: data <= 32'h00178793;         'd2187: data <= 32'h00f72023;
         'd2188: data <= 32'hfd1fe0ef;         'd2189: data <= 32'hf0091ce3;
         'd2190: data <= 32'hf11ff06f;         'd2191: data <= 32'h00090513;
         'd2192: data <= 32'h00c12083;         'd2193: data <= 32'h00812403;
         'd2194: data <= 32'h00412483;         'd2195: data <= 32'h00012903;
         'd2196: data <= 32'h01010113;         'd2197: data <= 32'h00008067;
         'd2198: data <= 32'h0a050663;         'd2199: data <= 32'hff010113;
         'd2200: data <= 32'h00112623;         'd2201: data <= 32'h00812423;
         'd2202: data <= 32'h00912223;         'd2203: data <= 32'h00050413;
         'd2204: data <= 32'hff050493;         'd2205: data <= 32'hff452783;
         'd2206: data <= 32'h0007c863;         'd2207: data <= 32'h30047073;
         'd2208: data <= 32'h00100073;         'd2209: data <= 32'h0000006f;
         'd2210: data <= 32'hff052703;         'd2211: data <= 32'h00070863;
         'd2212: data <= 32'h30047073;         'd2213: data <= 32'h00100073;
         'd2214: data <= 32'h0000006f;         'd2215: data <= 32'h0007cc63;
         'd2216: data <= 32'h00c12083;         'd2217: data <= 32'h00812403;
         'd2218: data <= 32'h00412483;         'd2219: data <= 32'h01010113;
         'd2220: data <= 32'h00008067;         'd2221: data <= 32'h80000737;
         'd2222: data <= 32'hfff74713;         'd2223: data <= 32'h00e7f7b3;
         'd2224: data <= 32'hfef52a23;         'd2225: data <= 32'hc8dfe0ef;
         'd2226: data <= 32'hff442683;         'd2227: data <= 32'h6fffe717;
         'd2228: data <= 32'hdb070713;         'd2229: data <= 32'h00072783;
         'd2230: data <= 32'h00d787b3;         'd2231: data <= 32'h00f72023;
         'd2232: data <= 32'h00048513;         'd2233: data <= 32'hd5dff0ef;
         'd2234: data <= 32'h6fffe717;         'd2235: data <= 32'hd8870713;
         'd2236: data <= 32'h00072783;         'd2237: data <= 32'h00178793;
         'd2238: data <= 32'h00f72023;         'd2239: data <= 32'hf05fe0ef;
         'd2240: data <= 32'hfa1ff06f;         'd2241: data <= 32'h00008067;
         'd2242: data <= 32'h00850793;         'd2243: data <= 32'h00f52223;
         'd2244: data <= 32'hfff00713;         'd2245: data <= 32'h00e52423;
         'd2246: data <= 32'h00f52623;         'd2247: data <= 32'h00f52823;
         'd2248: data <= 32'h00052023;         'd2249: data <= 32'h00008067;
         'd2250: data <= 32'h00052823;         'd2251: data <= 32'h00008067;
         'd2252: data <= 32'h0005a603;         'd2253: data <= 32'hfff00793;
         'd2254: data <= 32'h04f60063;         'd2255: data <= 32'h00850793;
         'd2256: data <= 32'h00078693;         'd2257: data <= 32'h0047a783;
         'd2258: data <= 32'h0007a703;         'd2259: data <= 32'hfee67ae3;
         'd2260: data <= 32'h0046a783;         'd2261: data <= 32'h00f5a223;
         'd2262: data <= 32'h00b7a423;         'd2263: data <= 32'h00d5a423;
         'd2264: data <= 32'h00b6a223;         'd2265: data <= 32'h00a5a823;
         'd2266: data <= 32'h00052783;         'd2267: data <= 32'h00178793;
         'd2268: data <= 32'h00f52023;         'd2269: data <= 32'h00008067;
         'd2270: data <= 32'h01052683;         'd2271: data <= 32'hfd5ff06f;
         'd2272: data <= 32'h01052783;         'd2273: data <= 32'h00452683;
         'd2274: data <= 32'h00852703;         'd2275: data <= 32'h00e6a423;
         'd2276: data <= 32'h00452683;         'd2277: data <= 32'h00d72223;
         'd2278: data <= 32'h0047a703;         'd2279: data <= 32'h00a70e63;
         'd2280: data <= 32'h00052823;         'd2281: data <= 32'h0007a703;
         'd2282: data <= 32'hfff70713;         'd2283: data <= 32'h00e7a023;
         'd2284: data <= 32'h0007a503;         'd2285: data <= 32'h00008067;
         'd2286: data <= 32'h00852703;         'd2287: data <= 32'h00e7a223;
         'd2288: data <= 32'hfe1ff06f;         'd2289: data <= 32'h30047073;
         'd2290: data <= 32'h6fffe717;         'd2291: data <= 32'hc4870713;
         'd2292: data <= 32'h00072783;         'd2293: data <= 32'h00178693;
         'd2294: data <= 32'h00d72023;         'd2295: data <= 32'h03852703;
         'd2296: data <= 32'h00071e63;         'd2297: data <= 32'h00100513;
         'd2298: data <= 32'h6fffe717;         'd2299: data <= 32'hc2f72423;
         'd2300: data <= 32'h00079463;         'd2301: data <= 32'h30046073;
         'd2302: data <= 32'h00008067;         'd2303: data <= 32'h00000513;
         'd2304: data <= 32'hfe9ff06f;         'd2305: data <= 32'h00050793;
         'd2306: data <= 32'h04052603;         'd2307: data <= 32'h04060063;
         'd2308: data <= 32'hff010113;         'd2309: data <= 32'h00112623;
         'd2310: data <= 32'h00058513;         'd2311: data <= 32'h00c7a703;
         'd2312: data <= 32'h00c70733;         'd2313: data <= 32'h00e7a623;
         'd2314: data <= 32'h0087a683;         'd2315: data <= 32'h00d76663;
         'd2316: data <= 32'h0007a703;         'd2317: data <= 32'h00e7a623;
         'd2318: data <= 32'h00c7a583;         'd2319: data <= 32'h7b0000ef;
         'd2320: data <= 32'h00c12083;         'd2321: data <= 32'h01010113;
         'd2322: data <= 32'h00008067;         'd2323: data <= 32'h00008067;
         'd2324: data <= 32'hff010113;         'd2325: data <= 32'h00112623;
         'd2326: data <= 32'h00812423;         'd2327: data <= 32'h00912223;
         'd2328: data <= 32'h00050493;         'd2329: data <= 32'h30047073;
         'd2330: data <= 32'h6fffe717;         'd2331: data <= 32'hba870713;
         'd2332: data <= 32'h00072783;         'd2333: data <= 32'h00178793;
         'd2334: data <= 32'h00f72023;         'd2335: data <= 32'h04554403;
         'd2336: data <= 32'h01841413;         'd2337: data <= 32'h41845413;
         'd2338: data <= 32'h0100006f;         'd2339: data <= 32'hfff40413;
         'd2340: data <= 32'h01841413;         'd2341: data <= 32'h41845413;
         'd2342: data <= 32'h02805063;         'd2343: data <= 32'h0244a783;
         'd2344: data <= 32'h00078c63;         'd2345: data <= 32'h02448513;
         'd2346: data <= 32'ha38ff0ef;         'd2347: data <= 32'hfe0500e3;
         'd2348: data <= 32'hce8ff0ef;         'd2349: data <= 32'hfd9ff06f;
         'd2350: data <= 32'hfff00793;         'd2351: data <= 32'h04f482a3;
         'd2352: data <= 32'h6fffe717;         'd2353: data <= 32'hb5070713;
         'd2354: data <= 32'h00072783;         'd2355: data <= 32'hfff78793;
         'd2356: data <= 32'h00f72023;         'd2357: data <= 32'h00079463;
         'd2358: data <= 32'h30046073;         'd2359: data <= 32'h30047073;
         'd2360: data <= 32'h6fffe717;         'd2361: data <= 32'hb3070713;
         'd2362: data <= 32'h00072783;         'd2363: data <= 32'h00178793;
         'd2364: data <= 32'h00f72023;         'd2365: data <= 32'h0444c403;
         'd2366: data <= 32'h01841413;         'd2367: data <= 32'h41845413;
         'd2368: data <= 32'h0100006f;         'd2369: data <= 32'hfff40413;
         'd2370: data <= 32'h01841413;         'd2371: data <= 32'h41845413;
         'd2372: data <= 32'h02805063;         'd2373: data <= 32'h0104a783;
         'd2374: data <= 32'h00078c63;         'd2375: data <= 32'h01048513;
         'd2376: data <= 32'h9c0ff0ef;         'd2377: data <= 32'hfe0500e3;
         'd2378: data <= 32'hc70ff0ef;         'd2379: data <= 32'hfd9ff06f;
         'd2380: data <= 32'hfff00793;         'd2381: data <= 32'h04f48223;
         'd2382: data <= 32'h6fffe717;         'd2383: data <= 32'had870713;
         'd2384: data <= 32'h00072783;         'd2385: data <= 32'hfff78793;
         'd2386: data <= 32'h00f72023;         'd2387: data <= 32'h00079463;
         'd2388: data <= 32'h30046073;         'd2389: data <= 32'h00c12083;
         'd2390: data <= 32'h00812403;         'd2391: data <= 32'h00412483;
         'd2392: data <= 32'h01010113;         'd2393: data <= 32'h00008067;
         'd2394: data <= 32'h10050c63;         'd2395: data <= 32'hfd010113;
         'd2396: data <= 32'h02112623;         'd2397: data <= 32'h02812423;
         'd2398: data <= 32'h02912223;         'd2399: data <= 32'h03212023;
         'd2400: data <= 32'h01312e23;         'd2401: data <= 32'h01412c23;
         'd2402: data <= 32'h01512a23;         'd2403: data <= 32'h01612823;
         'd2404: data <= 32'h01712623;         'd2405: data <= 32'h00050413;
         'd2406: data <= 32'h00058913;         'd2407: data <= 32'h03c52483;
         'd2408: data <= 32'h16048c63;         'd2409: data <= 32'h04052983;
         'd2410: data <= 32'h00000a13;         'd2411: data <= 32'h0104d693;
         'd2412: data <= 32'h0109d793;         'd2413: data <= 32'h12069263;
         'd2414: data <= 32'h01079713;         'd2415: data <= 32'h01075713;
         'd2416: data <= 32'h0c071663;         'd2417: data <= 32'h140a1a63;
         'd2418: data <= 32'h30047073;         'd2419: data <= 32'h6fffe717;
         'd2420: data <= 32'ha4470713;         'd2421: data <= 32'h00072783;
         'd2422: data <= 32'h00178793;         'd2423: data <= 32'h00f72023;
         'd2424: data <= 32'h00042483;         'd2425: data <= 32'h03c42a03;
         'd2426: data <= 32'h04042983;         'd2427: data <= 32'h00098593;
         'd2428: data <= 32'h000a0513;         'd2429: data <= 32'h0c5000ef;
         'd2430: data <= 32'h00a487b3;         'd2431: data <= 32'h00f42423;
         'd2432: data <= 32'h02042c23;         'd2433: data <= 32'h00942223;
         'd2434: data <= 32'hfffa0593;         'd2435: data <= 32'h00098513;
         'd2436: data <= 32'h0a9000ef;         'd2437: data <= 32'h00a484b3;
         'd2438: data <= 32'h00942623;         'd2439: data <= 32'hfff00793;
         'd2440: data <= 32'h04f40223;         'd2441: data <= 32'h04f402a3;
         'd2442: data <= 32'h0c091e63;         'd2443: data <= 32'h01042783;
         'd2444: data <= 32'h0c079063;         'd2445: data <= 32'h6fffe717;
         'd2446: data <= 32'h9dc70713;         'd2447: data <= 32'h00072783;
         'd2448: data <= 32'hfff78793;         'd2449: data <= 32'h00f72023;
         'd2450: data <= 32'h00079463;         'd2451: data <= 32'h30046073;
         'd2452: data <= 32'h00100513;         'd2453: data <= 32'h02c12083;
         'd2454: data <= 32'h02812403;         'd2455: data <= 32'h02412483;
         'd2456: data <= 32'h02012903;         'd2457: data <= 32'h01c12983;
         'd2458: data <= 32'h01812a03;         'd2459: data <= 32'h01412a83;
         'd2460: data <= 32'h01012b03;         'd2461: data <= 32'h00c12b83;
         'd2462: data <= 32'h03010113;         'd2463: data <= 32'h00008067;
         'd2464: data <= 32'h30047073;         'd2465: data <= 32'h00100073;
         'd2466: data <= 32'h0000006f;         'd2467: data <= 32'h00078b93;
         'd2468: data <= 32'h00048b13;         'd2469: data <= 32'h01099593;
         'd2470: data <= 32'h0105d593;         'd2471: data <= 32'h01049513;
         'd2472: data <= 32'h01055513;         'd2473: data <= 32'h015000ef;
         'd2474: data <= 32'h00050a93;         'd2475: data <= 32'h010b9593;
         'd2476: data <= 32'h0105d593;         'd2477: data <= 32'h010b1513;
         'd2478: data <= 32'h01055513;         'd2479: data <= 32'h7fc000ef;
         'd2480: data <= 32'h010ada93;         'd2481: data <= 32'h015507b3;
         'd2482: data <= 32'h0107d793;         'd2483: data <= 32'hee078ce3;
         'd2484: data <= 32'h00100a13;         'd2485: data <= 32'hef1ff06f;
         'd2486: data <= 32'h01079793;         'd2487: data <= 32'h0107d793;
         'd2488: data <= 32'hfe0798e3;         'd2489: data <= 32'h00068b93;
         'd2490: data <= 32'h00098b13;         'd2491: data <= 32'hfa9ff06f;
         'd2492: data <= 32'h01040513;         'd2493: data <= 32'hfedfe0ef;
         'd2494: data <= 32'hf2050ee3;         'd2495: data <= 32'h00000073;
         'd2496: data <= 32'hf35ff06f;         'd2497: data <= 32'h01040513;
         'd2498: data <= 32'hc01ff0ef;         'd2499: data <= 32'h02440513;
         'd2500: data <= 32'hbf9ff0ef;         'd2501: data <= 32'hf21ff06f;
         'd2502: data <= 32'h30047073;         'd2503: data <= 32'h00100073;
         'd2504: data <= 32'h0000006f;         'd2505: data <= 32'hff010113;
         'd2506: data <= 32'h00112623;         'd2507: data <= 32'h00050793;
         'd2508: data <= 32'h00070513;         'd2509: data <= 32'h02059263;
         'd2510: data <= 32'h00e52023;         'd2511: data <= 32'h02f52e23;
         'd2512: data <= 32'h04b52023;         'd2513: data <= 32'h00100593;
         'd2514: data <= 32'he21ff0ef;         'd2515: data <= 32'h00c12083;
         'd2516: data <= 32'h01010113;         'd2517: data <= 32'h00008067;
         'd2518: data <= 32'h00c72023;         'd2519: data <= 32'hfe1ff06f;
         'd2520: data <= 32'h12050663;         'd2521: data <= 32'hfe010113;
         'd2522: data <= 32'h00112e23;         'd2523: data <= 32'h00812c23;
         'd2524: data <= 32'h00912a23;         'd2525: data <= 32'h01212823;
         'd2526: data <= 32'h01312623;         'd2527: data <= 32'h01412423;
         'd2528: data <= 32'h01512223;         'd2529: data <= 32'h01612023;
         'd2530: data <= 32'h00050413;         'd2531: data <= 32'h00058493;
         'd2532: data <= 32'h00060913;         'd2533: data <= 32'h00000993;
         'd2534: data <= 32'h01055693;         'd2535: data <= 32'h0105d793;
         'd2536: data <= 32'h08069063;         'd2537: data <= 32'h01079713;
         'd2538: data <= 32'h01075713;         'd2539: data <= 32'h02071463;
         'd2540: data <= 32'h00099c63;         'd2541: data <= 32'h00048593;
         'd2542: data <= 32'h00040513;         'd2543: data <= 32'h6fc000ef;
         'd2544: data <= 32'hfb700793;         'd2545: data <= 32'h06a7fa63;
         'd2546: data <= 32'h30047073;         'd2547: data <= 32'h00100073;
         'd2548: data <= 32'h0000006f;         'd2549: data <= 32'h00078b13;
         'd2550: data <= 32'h00050a93;         'd2551: data <= 32'h01049593;
         'd2552: data <= 32'h0105d593;         'd2553: data <= 32'h01041513;
         'd2554: data <= 32'h01055513;         'd2555: data <= 32'h6cc000ef;
         'd2556: data <= 32'h00050a13;         'd2557: data <= 32'h010b1593;
         'd2558: data <= 32'h0105d593;         'd2559: data <= 32'h010a9513;
         'd2560: data <= 32'h01055513;         'd2561: data <= 32'h6b4000ef;
         'd2562: data <= 32'h010a5713;         'd2563: data <= 32'h00e507b3;
         'd2564: data <= 32'h0107d793;         'd2565: data <= 32'hf8078ee3;
         'd2566: data <= 32'h00100993;         'd2567: data <= 32'hf95ff06f;
         'd2568: data <= 32'h01079793;         'd2569: data <= 32'h0107d793;
         'd2570: data <= 32'hfe0798e3;         'd2571: data <= 32'h00068b13;
         'd2572: data <= 32'h00058a93;         'd2573: data <= 32'hfa9ff06f;
         'd2574: data <= 32'h04850513;         'd2575: data <= 32'h885ff0ef;
         'd2576: data <= 32'h00050993;         'd2577: data <= 32'h00050e63;
         'd2578: data <= 32'h00050713;         'd2579: data <= 32'h00090693;
         'd2580: data <= 32'h04850613;         'd2581: data <= 32'h00048593;
         'd2582: data <= 32'h00040513;         'd2583: data <= 32'hec9ff0ef;
         'd2584: data <= 32'h00098513;         'd2585: data <= 32'h01c12083;
         'd2586: data <= 32'h01812403;         'd2587: data <= 32'h01412483;
         'd2588: data <= 32'h01012903;         'd2589: data <= 32'h00c12983;
         'd2590: data <= 32'h00812a03;         'd2591: data <= 32'h00412a83;
         'd2592: data <= 32'h00012b03;         'd2593: data <= 32'h02010113;
         'd2594: data <= 32'h00008067;         'd2595: data <= 32'h30047073;
         'd2596: data <= 32'h00100073;         'd2597: data <= 32'h0000006f;
         'd2598: data <= 32'hfc010113;         'd2599: data <= 32'h02112e23;
         'd2600: data <= 32'h02812c23;         'd2601: data <= 32'h02912a23;
         'd2602: data <= 32'h03212823;         'd2603: data <= 32'h03312623;
         'd2604: data <= 32'h00c12623;         'd2605: data <= 32'h02050863;
         'd2606: data <= 32'h00050413;         'd2607: data <= 32'h00058913;
         'd2608: data <= 32'h02058863;         'd2609: data <= 32'h8e4ff0ef;
         'd2610: data <= 32'h00050493;         'd2611: data <= 32'h02051c63;
         'd2612: data <= 32'h00c12783;         'd2613: data <= 32'h10078263;
         'd2614: data <= 32'h30047073;         'd2615: data <= 32'h00100073;
         'd2616: data <= 32'h0000006f;         'd2617: data <= 32'h30047073;
         'd2618: data <= 32'h00100073;         'd2619: data <= 32'h0000006f;
         'd2620: data <= 32'h04052783;         'd2621: data <= 32'hfc0788e3;
         'd2622: data <= 32'h30047073;         'd2623: data <= 32'h00100073;
         'd2624: data <= 32'h0000006f;         'd2625: data <= 32'h00000493;
         'd2626: data <= 32'h0d00006f;         'd2627: data <= 32'h00090593;
         'd2628: data <= 32'h00040513;         'd2629: data <= 32'haf1ff0ef;
         'd2630: data <= 32'hfff98993;         'd2631: data <= 32'h03342c23;
         'd2632: data <= 32'h01042783;         'd2633: data <= 32'h04079063;
         'd2634: data <= 32'h6fffd717;         'd2635: data <= 32'h6e870713;
         'd2636: data <= 32'h00072783;         'd2637: data <= 32'hfff78793;
         'd2638: data <= 32'h00f72023;         'd2639: data <= 32'h00079463;
         'd2640: data <= 32'h30046073;         'd2641: data <= 32'h00100513;
         'd2642: data <= 32'h03c12083;         'd2643: data <= 32'h03812403;
         'd2644: data <= 32'h03412483;         'd2645: data <= 32'h03012903;
         'd2646: data <= 32'h02c12983;         'd2647: data <= 32'h04010113;
         'd2648: data <= 32'h00008067;         'd2649: data <= 32'h01040513;
         'd2650: data <= 32'hd79fe0ef;         'd2651: data <= 32'hfa050ee3;
         'd2652: data <= 32'h00000073;         'd2653: data <= 32'hfb5ff06f;
         'd2654: data <= 32'h6fffd797;         'd2655: data <= 32'h68e7ac23;
         'd2656: data <= 32'h00071463;         'd2657: data <= 32'h30046073;
         'd2658: data <= 32'h00000513;         'd2659: data <= 32'hfbdff06f;
         'd2660: data <= 32'h01810513;         'd2661: data <= 32'hed5fe0ef;
         'd2662: data <= 32'h00100493;         'd2663: data <= 32'h0680006f;
         'd2664: data <= 32'h04040223;         'd2665: data <= 32'h0ac0006f;
         'd2666: data <= 32'h040402a3;         'd2667: data <= 32'h0b80006f;
         'd2668: data <= 32'h00040513;         'd2669: data <= 32'ha9dff0ef;
         'd2670: data <= 32'h849fe0ef;         'd2671: data <= 32'h01c0006f;
         'd2672: data <= 32'h00040513;         'd2673: data <= 32'ha8dff0ef;
         'd2674: data <= 32'h839fe0ef;         'd2675: data <= 32'h00040513;
         'd2676: data <= 32'h9f5ff0ef;         'd2677: data <= 32'h0e051063;
         'd2678: data <= 32'h30047073;         'd2679: data <= 32'h6fffd797;
         'd2680: data <= 32'h63478793;         'd2681: data <= 32'h0007a703;
         'd2682: data <= 32'h00170693;         'd2683: data <= 32'h00d7a023;
         'd2684: data <= 32'h03842983;         'd2685: data <= 32'hf0099ce3;
         'd2686: data <= 32'h00c12783;         'd2687: data <= 32'hf6078ee3;
         'd2688: data <= 32'hf80488e3;         'd2689: data <= 32'h6fffd717;
         'd2690: data <= 32'h60c70713;         'd2691: data <= 32'h00072783;
         'd2692: data <= 32'hfff78793;         'd2693: data <= 32'h00f72023;
         'd2694: data <= 32'h00079463;         'd2695: data <= 32'h30046073;
         'd2696: data <= 32'hd30fe0ef;         'd2697: data <= 32'h30047073;
         'd2698: data <= 32'h6fffd717;         'd2699: data <= 32'h5e870713;
         'd2700: data <= 32'h00072783;         'd2701: data <= 32'h00178693;
         'd2702: data <= 32'h00d72023;         'd2703: data <= 32'h04444703;
         'd2704: data <= 32'h01871713;         'd2705: data <= 32'h41875713;
         'd2706: data <= 32'hfff00693;         'd2707: data <= 32'hf4d70ae3;
         'd2708: data <= 32'h04544703;         'd2709: data <= 32'h01871713;
         'd2710: data <= 32'h41875713;         'd2711: data <= 32'hfff00693;
         'd2712: data <= 32'hf4d704e3;         'd2713: data <= 32'h6fffd717;
         'd2714: data <= 32'h5af72623;         'd2715: data <= 32'h00079463;
         'd2716: data <= 32'h30046073;         'd2717: data <= 32'h00c10593;
         'd2718: data <= 32'h01810513;         'd2719: data <= 32'he09fe0ef;
         'd2720: data <= 32'hf40510e3;         'd2721: data <= 32'h00040513;
         'd2722: data <= 32'h93dff0ef;         'd2723: data <= 32'hf20502e3;
         'd2724: data <= 32'h00c12583;         'd2725: data <= 32'h02440513;
         'd2726: data <= 32'hb75fe0ef;         'd2727: data <= 32'h00040513;
         'd2728: data <= 32'h9b1ff0ef;         'd2729: data <= 32'hf5cfe0ef;
         'd2730: data <= 32'hf20518e3;         'd2731: data <= 32'h00000073;
         'd2732: data <= 32'hf29ff06f;         'd2733: data <= 32'h00000513;
         'd2734: data <= 32'he91ff06f;         'd2735: data <= 32'h00050a63;
         'd2736: data <= 32'h00058e63;         'd2737: data <= 32'h00000613;
         'd2738: data <= 32'h00000793;         'd2739: data <= 32'h0280006f;
         'd2740: data <= 32'h30047073;         'd2741: data <= 32'h00100073;
         'd2742: data <= 32'h0000006f;         'd2743: data <= 32'h00008067;
         'd2744: data <= 32'h6ffff617;         'd2745: data <= 32'h2b060613;
         'd2746: data <= 32'h00c68633;         'd2747: data <= 32'h0580006f;
         'd2748: data <= 32'h00178793;         'd2749: data <= 32'h00700713;
         'd2750: data <= 32'h04f76463;         'd2751: data <= 32'h00379693;
         'd2752: data <= 32'h6ffff717;         'd2753: data <= 32'h29070713;
         'd2754: data <= 32'h00d70733;         'd2755: data <= 32'h00472703;
         'd2756: data <= 32'hfca708e3;         'd2757: data <= 32'hfc061ee3;
         'd2758: data <= 32'h00379693;         'd2759: data <= 32'h6ffff717;
         'd2760: data <= 32'h27470713;         'd2761: data <= 32'h00d70733;
         'd2762: data <= 32'h00072703;         'd2763: data <= 32'hfc0712e3;
         'd2764: data <= 32'h6ffff717;         'd2765: data <= 32'h26070713;
         'd2766: data <= 32'h00e68633;         'd2767: data <= 32'hfb5ff06f;
         'd2768: data <= 32'h00060663;         'd2769: data <= 32'h00b62023;
         'd2770: data <= 32'h00a62223;         'd2771: data <= 32'h00008067;
         'd2772: data <= 32'hff010113;         'd2773: data <= 32'h00112623;
         'd2774: data <= 32'h00812423;         'd2775: data <= 32'h00050413;
         'd2776: data <= 32'h30047073;         'd2777: data <= 32'h6fffd717;
         'd2778: data <= 32'h4ac70713;         'd2779: data <= 32'h00072783;
         'd2780: data <= 32'h00178693;         'd2781: data <= 32'h00d72023;
         'd2782: data <= 32'h04454703;         'd2783: data <= 32'h01871713;
         'd2784: data <= 32'h41875713;         'd2785: data <= 32'hfff00693;
         'd2786: data <= 32'h04d70463;         'd2787: data <= 32'h04544703;
         'd2788: data <= 32'h01871713;         'd2789: data <= 32'h41875713;
         'd2790: data <= 32'hfff00693;         'd2791: data <= 32'h02d70e63;
         'd2792: data <= 32'h6fffd717;         'd2793: data <= 32'h46f72823;
         'd2794: data <= 32'h00079463;         'd2795: data <= 32'h30046073;
         'd2796: data <= 32'h03842783;         'd2797: data <= 32'h02078663;
         'd2798: data <= 32'h00040513;         'd2799: data <= 32'h895ff0ef;
         'd2800: data <= 32'h00c12083;         'd2801: data <= 32'h00812403;
         'd2802: data <= 32'h01010113;         'd2803: data <= 32'h00008067;
         'd2804: data <= 32'h04050223;         'd2805: data <= 32'hfb9ff06f;
         'd2806: data <= 32'h040402a3;         'd2807: data <= 32'hfc5ff06f;
         'd2808: data <= 32'h02440513;         'd2809: data <= 32'ha75fe0ef;
         'd2810: data <= 32'hfd1ff06f;         'd2811: data <= 32'h00b547b3;
         'd2812: data <= 32'h0037f793;         'd2813: data <= 32'h00c508b3;
         'd2814: data <= 32'h06079463;         'd2815: data <= 32'h00300793;
         'd2816: data <= 32'h06c7f063;         'd2817: data <= 32'h00357793;
         'd2818: data <= 32'h00050713;         'd2819: data <= 32'h06079a63;
         'd2820: data <= 32'hffc8f613;         'd2821: data <= 32'h40e606b3;
         'd2822: data <= 32'h02000793;         'd2823: data <= 32'h08d7ce63;
         'd2824: data <= 32'h00058693;         'd2825: data <= 32'h00070793;
         'd2826: data <= 32'h02c77863;         'd2827: data <= 32'h0006a803;
         'd2828: data <= 32'h00478793;         'd2829: data <= 32'h00468693;
         'd2830: data <= 32'hff07ae23;         'd2831: data <= 32'hfec7e8e3;
         'd2832: data <= 32'hfff60793;         'd2833: data <= 32'h40e787b3;
         'd2834: data <= 32'hffc7f793;         'd2835: data <= 32'h00478793;
         'd2836: data <= 32'h00f70733;         'd2837: data <= 32'h00f585b3;
         'd2838: data <= 32'h01176863;         'd2839: data <= 32'h00008067;
         'd2840: data <= 32'h00050713;         'd2841: data <= 32'h05157863;
         'd2842: data <= 32'h0005c783;         'd2843: data <= 32'h00170713;
         'd2844: data <= 32'h00158593;         'd2845: data <= 32'hfef70fa3;
         'd2846: data <= 32'hfee898e3;         'd2847: data <= 32'h00008067;
         'd2848: data <= 32'h0005c683;         'd2849: data <= 32'h00170713;
         'd2850: data <= 32'h00377793;         'd2851: data <= 32'hfed70fa3;
         'd2852: data <= 32'h00158593;         'd2853: data <= 32'hf6078ee3;
         'd2854: data <= 32'h0005c683;         'd2855: data <= 32'h00170713;
         'd2856: data <= 32'h00377793;         'd2857: data <= 32'hfed70fa3;
         'd2858: data <= 32'h00158593;         'd2859: data <= 32'hfc079ae3;
         'd2860: data <= 32'hf61ff06f;         'd2861: data <= 32'h00008067;
         'd2862: data <= 32'hff010113;         'd2863: data <= 32'h00812623;
         'd2864: data <= 32'h02000413;         'd2865: data <= 32'h0005a383;
         'd2866: data <= 32'h0045a283;         'd2867: data <= 32'h0085af83;
         'd2868: data <= 32'h00c5af03;         'd2869: data <= 32'h0105ae83;
         'd2870: data <= 32'h0145ae03;         'd2871: data <= 32'h0185a303;
         'd2872: data <= 32'h01c5a803;         'd2873: data <= 32'h0205a683;
         'd2874: data <= 32'h02470713;         'd2875: data <= 32'h40e607b3;
         'd2876: data <= 32'hfc772e23;         'd2877: data <= 32'hfe572023;
         'd2878: data <= 32'hfff72223;         'd2879: data <= 32'hffe72423;
         'd2880: data <= 32'hffd72623;         'd2881: data <= 32'hffc72823;
         'd2882: data <= 32'hfe672a23;         'd2883: data <= 32'hff072c23;
         'd2884: data <= 32'hfed72e23;         'd2885: data <= 32'h02458593;
         'd2886: data <= 32'hfaf446e3;         'd2887: data <= 32'h00058693;
         'd2888: data <= 32'h00070793;         'd2889: data <= 32'h02c77863;
         'd2890: data <= 32'h0006a803;         'd2891: data <= 32'h00478793;
         'd2892: data <= 32'h00468693;         'd2893: data <= 32'hff07ae23;
         'd2894: data <= 32'hfec7e8e3;         'd2895: data <= 32'hfff60793;
         'd2896: data <= 32'h40e787b3;         'd2897: data <= 32'hffc7f793;
         'd2898: data <= 32'h00478793;         'd2899: data <= 32'h00f70733;
         'd2900: data <= 32'h00f585b3;         'd2901: data <= 32'h01176863;
         'd2902: data <= 32'h00c12403;         'd2903: data <= 32'h01010113;
         'd2904: data <= 32'h00008067;         'd2905: data <= 32'h0005c783;
         'd2906: data <= 32'h00170713;         'd2907: data <= 32'h00158593;
         'd2908: data <= 32'hfef70fa3;         'd2909: data <= 32'hfee882e3;
         'd2910: data <= 32'h0005c783;         'd2911: data <= 32'h00170713;
         'd2912: data <= 32'h00158593;         'd2913: data <= 32'hfef70fa3;
         'd2914: data <= 32'hfce89ee3;         'd2915: data <= 32'hfcdff06f;
         'd2916: data <= 32'h00f00313;         'd2917: data <= 32'h00050713;
         'd2918: data <= 32'h02c37e63;         'd2919: data <= 32'h00f77793;
         'd2920: data <= 32'h0a079063;         'd2921: data <= 32'h08059263;
         'd2922: data <= 32'hff067693;         'd2923: data <= 32'h00f67613;
         'd2924: data <= 32'h00e686b3;         'd2925: data <= 32'h00b72023;
         'd2926: data <= 32'h00b72223;         'd2927: data <= 32'h00b72423;
         'd2928: data <= 32'h00b72623;         'd2929: data <= 32'h01070713;
         'd2930: data <= 32'hfed766e3;         'd2931: data <= 32'h00061463;
         'd2932: data <= 32'h00008067;         'd2933: data <= 32'h40c306b3;
         'd2934: data <= 32'h00269693;         'd2935: data <= 32'h00000297;
         'd2936: data <= 32'h005686b3;         'd2937: data <= 32'h00c68067;
         'd2938: data <= 32'h00b70723;         'd2939: data <= 32'h00b706a3;
         'd2940: data <= 32'h00b70623;         'd2941: data <= 32'h00b705a3;
         'd2942: data <= 32'h00b70523;         'd2943: data <= 32'h00b704a3;
         'd2944: data <= 32'h00b70423;         'd2945: data <= 32'h00b703a3;
         'd2946: data <= 32'h00b70323;         'd2947: data <= 32'h00b702a3;
         'd2948: data <= 32'h00b70223;         'd2949: data <= 32'h00b701a3;
         'd2950: data <= 32'h00b70123;         'd2951: data <= 32'h00b700a3;
         'd2952: data <= 32'h00b70023;         'd2953: data <= 32'h00008067;
         'd2954: data <= 32'h0ff5f593;         'd2955: data <= 32'h00859693;
         'd2956: data <= 32'h00d5e5b3;         'd2957: data <= 32'h01059693;
         'd2958: data <= 32'h00d5e5b3;         'd2959: data <= 32'hf6dff06f;
         'd2960: data <= 32'h00279693;         'd2961: data <= 32'h00000297;
         'd2962: data <= 32'h005686b3;         'd2963: data <= 32'h00008293;
         'd2964: data <= 32'hfa0680e7;         'd2965: data <= 32'h00028093;
         'd2966: data <= 32'hff078793;         'd2967: data <= 32'h40f70733;
         'd2968: data <= 32'h00f60633;         'd2969: data <= 32'hf6c378e3;
         'd2970: data <= 32'hf3dff06f;         'd2971: data <= 32'h000107b7;
         'd2972: data <= 32'h02f57a63;         'd2973: data <= 32'h10053793;
         'd2974: data <= 32'h0017c793;         'd2975: data <= 32'h00379793;
         'd2976: data <= 32'ha0003737;         'd2977: data <= 32'h02000693;
         'd2978: data <= 32'h40f686b3;         'd2979: data <= 32'h00f55533;
         'd2980: data <= 32'h65870793;         'd2981: data <= 32'h00a787b3;
         'd2982: data <= 32'h0007c503;         'd2983: data <= 32'h40a68533;
         'd2984: data <= 32'h00008067;         'd2985: data <= 32'h01000737;
         'd2986: data <= 32'h01000793;         'd2987: data <= 32'hfce56ae3;
         'd2988: data <= 32'h01800793;         'd2989: data <= 32'hfcdff06f;
         'd2990: data <= 32'h00050613;         'd2991: data <= 32'h00000513;
         'd2992: data <= 32'h0015f693;         'd2993: data <= 32'h00068463;
         'd2994: data <= 32'h00c50533;         'd2995: data <= 32'h0015d593;
         'd2996: data <= 32'h00161613;         'd2997: data <= 32'hfe0596e3;
         'd2998: data <= 32'h00008067;         'd2999: data <= 32'h06054063;
         'd3000: data <= 32'h0605c663;         'd3001: data <= 32'h00058613;
         'd3002: data <= 32'h00050593;         'd3003: data <= 32'hfff00513;
         'd3004: data <= 32'h02060c63;         'd3005: data <= 32'h00100693;
         'd3006: data <= 32'h00b67a63;         'd3007: data <= 32'h00c05863;
         'd3008: data <= 32'h00161613;         'd3009: data <= 32'h00169693;
         'd3010: data <= 32'hfeb66ae3;         'd3011: data <= 32'h00000513;
         'd3012: data <= 32'h00c5e663;         'd3013: data <= 32'h40c585b3;
         'd3014: data <= 32'h00d56533;         'd3015: data <= 32'h0016d693;
         'd3016: data <= 32'h00165613;         'd3017: data <= 32'hfe0696e3;
         'd3018: data <= 32'h00008067;         'd3019: data <= 32'h00008293;
         'd3020: data <= 32'hfb5ff0ef;         'd3021: data <= 32'h00058513;
         'd3022: data <= 32'h00028067;         'd3023: data <= 32'h40a00533;
         'd3024: data <= 32'h00b04863;         'd3025: data <= 32'h40b005b3;
         'd3026: data <= 32'hf9dff06f;         'd3027: data <= 32'h40b005b3;
         'd3028: data <= 32'h00008293;         'd3029: data <= 32'hf91ff0ef;
         'd3030: data <= 32'h40a00533;         'd3031: data <= 32'h00028067;
         'd3032: data <= 32'h00008293;         'd3033: data <= 32'h0005ca63;
         'd3034: data <= 32'h00054c63;         'd3035: data <= 32'hf79ff0ef;
         'd3036: data <= 32'h00058513;         'd3037: data <= 32'h00028067;
         'd3038: data <= 32'h40b005b3;         'd3039: data <= 32'hfe0558e3;
         'd3040: data <= 32'h40a00533;         'd3041: data <= 32'hf61ff0ef;
         'd3042: data <= 32'h40b00533;         'd3043: data <= 32'h00028067;
         'd3044: data <= 32'hff010113;         'd3045: data <= 32'hf14027f3;
         'd3046: data <= 32'h00f12623;         'd3047: data <= 32'h00c12603;
         'd3048: data <= 32'h1e0007b7;         'd3049: data <= 32'h00178793;
         'd3050: data <= 32'h00f60633;         'd3051: data <= 32'h00361613;
         'd3052: data <= 32'h6fffd797;         'd3053: data <= 32'h0ec7a023;
         'd3054: data <= 32'hf00007b7;         'd3055: data <= 32'h0047a703;
         'd3056: data <= 32'h0007a683;         'd3057: data <= 32'h0047a783;
         'd3058: data <= 32'hfee798e3;         'd3059: data <= 32'h6fffd797;
         'd3060: data <= 32'h0cc78793;         'd3061: data <= 32'h00e7a023;
         'd3062: data <= 32'h0007a223;         'd3063: data <= 32'h0007a023;
         'd3064: data <= 32'h00e7a223;         'd3065: data <= 32'h00d7a023;
         'd3066: data <= 32'h000185b7;         'd3067: data <= 32'h6a058593;
         'd3068: data <= 32'h00b685b3;         'd3069: data <= 32'h00d5b533;
         'd3070: data <= 32'h00e508b3;         'd3071: data <= 32'h00b7a023;
         'd3072: data <= 32'h0117a223;         'd3073: data <= 32'h00b62023;
         'd3074: data <= 32'h01162223;         'd3075: data <= 32'h00031637;
         'd3076: data <= 32'hd4060613;         'd3077: data <= 32'h00c68633;
         'd3078: data <= 32'h00d636b3;         'd3079: data <= 32'h00e686b3;
         'd3080: data <= 32'h00c7a023;         'd3081: data <= 32'h00d7a223;
         'd3082: data <= 32'h01010113;         'd3083: data <= 32'h00008067;
         'd3084: data <= 32'hff010113;         'd3085: data <= 32'h00112623;
         'd3086: data <= 32'h20000613;         'd3087: data <= 32'h0ee00593;
         'd3088: data <= 32'h6ffff517;         'd3089: data <= 32'hd9050513;
         'd3090: data <= 32'hd49ff0ef;         'd3091: data <= 32'hf45ff0ef;
         'd3092: data <= 32'h000017b7;         'd3093: data <= 32'h88078793;
         'd3094: data <= 32'h3047a073;         'd3095: data <= 32'h074000ef;
         'd3096: data <= 32'h00000513;         'd3097: data <= 32'h00c12083;
         'd3098: data <= 32'h01010113;         'd3099: data <= 32'h00008067;
         'd3100: data <= 32'h300022f3;         'd3101: data <= 32'hff72f293;
         'd3102: data <= 32'h18800313;         'd3103: data <= 32'h00431313;
         'd3104: data <= 32'h0062e2b3;         'd3105: data <= 32'hffc50513;
         'd3106: data <= 32'h00552023;         'd3107: data <= 32'hffc50513;
         'd3108: data <= 32'h00052023;         'd3109: data <= 32'hfa850513;
         'd3110: data <= 32'h00c52023;         'd3111: data <= 32'hfe850513;
         'd3112: data <= 32'h6fffd297;         'd3113: data <= 32'hfec2a283;
         'd3114: data <= 32'h00552023;         'd3115: data <= 32'h00000293;
         'd3116: data <= 32'h00028a63;         'd3117: data <= 32'hffc50513;
         'd3118: data <= 32'h00052023;         'd3119: data <= 32'hfff28293;
         'd3120: data <= 32'hff1ff06f;         'd3121: data <= 32'hffc50513;
         'd3122: data <= 32'h00b52023;         'd3123: data <= 32'h00008067;
         'd3124: data <= 32'h6fffd117;         'd3125: data <= 32'hf8812103;
         'd3126: data <= 32'h00012103;         'd3127: data <= 32'h00012083;
         'd3128: data <= 32'h01012383;         'd3129: data <= 32'h01412403;
         'd3130: data <= 32'h01812483;         'd3131: data <= 32'h01c12503;
         'd3132: data <= 32'h02012583;         'd3133: data <= 32'h02412603;
         'd3134: data <= 32'h02812683;         'd3135: data <= 32'h02c12703;
         'd3136: data <= 32'h03012783;         'd3137: data <= 32'h03412803;
         'd3138: data <= 32'h03812883;         'd3139: data <= 32'h03c12903;
         'd3140: data <= 32'h04012983;         'd3141: data <= 32'h04412a03;
         'd3142: data <= 32'h04812a83;         'd3143: data <= 32'h04c12b03;
         'd3144: data <= 32'h05012b83;         'd3145: data <= 32'h05412c03;
         'd3146: data <= 32'h05812c83;         'd3147: data <= 32'h05c12d03;
         'd3148: data <= 32'h06012d83;         'd3149: data <= 32'h06412e03;
         'd3150: data <= 32'h06812e83;         'd3151: data <= 32'h06c12f03;
         'd3152: data <= 32'h07012f83;         'd3153: data <= 32'h07412283;
         'd3154: data <= 32'h6fffd317;         'd3155: data <= 32'hec432303;
         'd3156: data <= 32'h00532023;         'd3157: data <= 32'h07812283;
         'd3158: data <= 32'h00828293;         'd3159: data <= 32'h30029073;
         'd3160: data <= 32'h00812283;         'd3161: data <= 32'h00c12303;
         'd3162: data <= 32'h07c10113;         'd3163: data <= 32'h00008067;
         'd3164: data <= 32'h342022f3;         'd3165: data <= 32'h34102373;
         'd3166: data <= 32'h300023f3;         'd3167: data <= 32'h0000006f;
         'd3168: data <= 32'h342022f3;         'd3169: data <= 32'h34102373;
         'd3170: data <= 32'h300023f3;         'd3171: data <= 32'h0000006f;
         'd3172: data <= 32'h00000000;         'd3173: data <= 32'h00000000;
         'd3174: data <= 32'h00000000;         'd3175: data <= 32'h00000000;
         'd3176: data <= 32'h00000000;         'd3177: data <= 32'h00000000;
         'd3178: data <= 32'h00000000;         'd3179: data <= 32'h00000000;
         'd3180: data <= 32'h00000000;         'd3181: data <= 32'h00000000;
         'd3182: data <= 32'h00000000;         'd3183: data <= 32'h00000000;
         'd3184: data <= 32'h00000000;         'd3185: data <= 32'h00000000;
         'd3186: data <= 32'h00000000;         'd3187: data <= 32'h00000000;
         'd3188: data <= 32'h00000000;         'd3189: data <= 32'h00000000;
         'd3190: data <= 32'h00000000;         'd3191: data <= 32'h00000000;
         'd3192: data <= 32'h00000000;         'd3193: data <= 32'h00000000;
         'd3194: data <= 32'h00000000;         'd3195: data <= 32'h00000000;
         'd3196: data <= 32'h00000000;         'd3197: data <= 32'h00000000;
         'd3198: data <= 32'h00000000;         'd3199: data <= 32'h00000000;
         'd3200: data <= 32'hf8410113;         'd3201: data <= 32'h00112223;
         'd3202: data <= 32'h00512423;         'd3203: data <= 32'h00612623;
         'd3204: data <= 32'h00712823;         'd3205: data <= 32'h00812a23;
         'd3206: data <= 32'h00912c23;         'd3207: data <= 32'h00a12e23;
         'd3208: data <= 32'h02b12023;         'd3209: data <= 32'h02c12223;
         'd3210: data <= 32'h02d12423;         'd3211: data <= 32'h02e12623;
         'd3212: data <= 32'h02f12823;         'd3213: data <= 32'h03012a23;
         'd3214: data <= 32'h03112c23;         'd3215: data <= 32'h03212e23;
         'd3216: data <= 32'h05312023;         'd3217: data <= 32'h05412223;
         'd3218: data <= 32'h05512423;         'd3219: data <= 32'h05612623;
         'd3220: data <= 32'h05712823;         'd3221: data <= 32'h05812a23;
         'd3222: data <= 32'h05912c23;         'd3223: data <= 32'h05a12e23;
         'd3224: data <= 32'h07b12023;         'd3225: data <= 32'h07c12223;
         'd3226: data <= 32'h07d12423;         'd3227: data <= 32'h07e12623;
         'd3228: data <= 32'h07f12823;         'd3229: data <= 32'h6fffd297;
         'd3230: data <= 32'hd9c2a283;         'd3231: data <= 32'h06512a23;
         'd3232: data <= 32'h300022f3;         'd3233: data <= 32'h06512c23;
         'd3234: data <= 32'h6fffd297;         'd3235: data <= 32'hdd02a283;
         'd3236: data <= 32'h0022a023;         'd3237: data <= 32'h34202573;
         'd3238: data <= 32'h341025f3;         'd3239: data <= 32'h00055a63;
         'd3240: data <= 32'h00b12023;         'd3241: data <= 32'h6fffd117;
         'd3242: data <= 32'hd6012103;         'd3243: data <= 32'h0180006f;
         'd3244: data <= 32'h00458593;         'd3245: data <= 32'h00b12023;
         'd3246: data <= 32'h6fffd117;         'd3247: data <= 32'hd4c12103;
         'd3248: data <= 32'h0700006f;         'd3249: data <= 32'h00100293;
         'd3250: data <= 32'h01f29293;         'd3251: data <= 32'h00728313;
         'd3252: data <= 32'h04651c63;         'd3253: data <= 32'h6fffd517;
         'd3254: data <= 32'hdbc52503;         'd3255: data <= 32'h6fffd597;
         'd3256: data <= 32'hd385a583;         'd3257: data <= 32'hfff00713;
         'd3258: data <= 32'h0005a603;         'd3259: data <= 32'h0045a683;
         'd3260: data <= 32'h00e52023;         'd3261: data <= 32'h00d52223;
         'd3262: data <= 32'h00c52023;         'd3263: data <= 32'h6fffd297;
         'd3264: data <= 32'hd042a283;         'd3265: data <= 32'h00c28733;
         'd3266: data <= 32'h00c73333;         'd3267: data <= 32'h006683b3;
         'd3268: data <= 32'h00e5a023;         'd3269: data <= 32'h0075a223;
         'd3270: data <= 32'hc5dfd0ef;         'd3271: data <= 32'h02050663;
         'd3272: data <= 32'h994fe0ef;         'd3273: data <= 32'h0240006f;
         'd3274: data <= 32'h83cfd0ef;         'd3275: data <= 32'h01c0006f;
         'd3276: data <= 32'h00b00293;         'd3277: data <= 32'h00551663;
         'd3278: data <= 32'h97cfe0ef;         'd3279: data <= 32'h00c0006f;
         'd3280: data <= 32'h868fd0ef;         'd3281: data <= 32'h0040006f;
         'd3282: data <= 32'h6fffd317;         'd3283: data <= 32'hd1032303;
         'd3284: data <= 32'h00032103;         'd3285: data <= 32'h00012283;
         'd3286: data <= 32'h34129073;         'd3287: data <= 32'h07812283;
         'd3288: data <= 32'h30029073;         'd3289: data <= 32'h07412283;
         'd3290: data <= 32'h6fffd317;         'd3291: data <= 32'hca432303;
         'd3292: data <= 32'h00532023;         'd3293: data <= 32'h00412083;
         'd3294: data <= 32'h00812283;         'd3295: data <= 32'h00c12303;
         'd3296: data <= 32'h01012383;         'd3297: data <= 32'h01412403;
         'd3298: data <= 32'h01812483;         'd3299: data <= 32'h01c12503;
         'd3300: data <= 32'h02012583;         'd3301: data <= 32'h02412603;
         'd3302: data <= 32'h02812683;         'd3303: data <= 32'h02c12703;
         'd3304: data <= 32'h03012783;         'd3305: data <= 32'h03412803;
         'd3306: data <= 32'h03812883;         'd3307: data <= 32'h03c12903;
         'd3308: data <= 32'h04012983;         'd3309: data <= 32'h04412a03;
         'd3310: data <= 32'h04812a83;         'd3311: data <= 32'h04c12b03;
         'd3312: data <= 32'h05012b83;         'd3313: data <= 32'h05412c03;
         'd3314: data <= 32'h05812c83;         'd3315: data <= 32'h05c12d03;
         'd3316: data <= 32'h06012d83;         'd3317: data <= 32'h06412e03;
         'd3318: data <= 32'h06812e83;         'd3319: data <= 32'h06c12f03;
         'd3320: data <= 32'h07012f83;         'd3321: data <= 32'h07c10113;
         'd3322: data <= 32'h30200073;         'd3323: data <= 32'h00000000;
         'd3324: data <= 32'h7361540a;         'd3325: data <= 32'h202d206b;
         'd3326: data <= 32'h202f2034;         'd3327: data <= 32'h74736554;
         'd3328: data <= 32'h6425203a;         'd3329: data <= 32'h00000000;
         'd3330: data <= 32'h7361540a;         'd3331: data <= 32'h202d206b;
         'd3332: data <= 32'h202f2033;         'd3333: data <= 32'h74736554;
         'd3334: data <= 32'h6425203a;         'd3335: data <= 32'h00000000;
         'd3336: data <= 32'h7361540a;         'd3337: data <= 32'h202d206b;
         'd3338: data <= 32'h202f2032;         'd3339: data <= 32'h74736554;
         'd3340: data <= 32'h6425203a;         'd3341: data <= 32'h00000000;
         'd3342: data <= 32'h7361540a;         'd3343: data <= 32'h202d206b;
         'd3344: data <= 32'h202f2031;         'd3345: data <= 32'h74736554;
         'd3346: data <= 32'h6425203a;         'd3347: data <= 32'h00000000;
         'd3348: data <= 32'h00003154;         'd3349: data <= 32'h00003249;
         'd3350: data <= 32'h00003354;         'd3351: data <= 32'h00003454;
         'd3352: data <= 32'h2e303156;         'd3353: data <= 32'h2b342e34;
         'd3354: data <= 32'h00000000;         'd3355: data <= 32'h6572460a;
         'd3356: data <= 32'h4f545265;         'd3357: data <= 32'h73252053;
         'd3358: data <= 32'h206e6f20;         'd3359: data <= 32'h20586f4e;
         'd3360: data <= 32'h20436f53;         'd3361: data <= 32'h6f6d6544;
         'd3362: data <= 32'h00000a0a;         'd3363: data <= 32'h0a63250a;
         'd3364: data <= 32'h00000000;         'd3365: data <= 32'h52493c0a;
         'd3366: data <= 32'h6d203e51;         'd3367: data <= 32'h73756163;
         'd3368: data <= 32'h203d2065;         'd3369: data <= 32'h78257830;
         'd3370: data <= 32'h492f3c20;         'd3371: data <= 32'h0a3e5152;
         'd3372: data <= 32'h00000000;         'd3373: data <= 32'h58453c0a;
         'd3374: data <= 32'h6d203e43;         'd3375: data <= 32'h73756163;
         'd3376: data <= 32'h203d2065;         'd3377: data <= 32'h78257830;
         'd3378: data <= 32'h452f3c20;         'd3379: data <= 32'h0a3e4358;
         'd3380: data <= 32'h00000000;         'd3381: data <= 32'h65657246;
         'd3382: data <= 32'h534f5452;         'd3383: data <= 32'h5541465f;
         'd3384: data <= 32'h203a544c;         'd3385: data <= 32'h70704176;
         'd3386: data <= 32'h6163696c;         'd3387: data <= 32'h6e6f6974;
         'd3388: data <= 32'h6c6c614d;         'd3389: data <= 32'h6146636f;
         'd3390: data <= 32'h64656c69;         'd3391: data <= 32'h6b6f6f48;
         'd3392: data <= 32'h6f732820;         'd3393: data <= 32'h6974756c;
         'd3394: data <= 32'h203a6e6f;         'd3395: data <= 32'h72636e69;
         'd3396: data <= 32'h65736165;         'd3397: data <= 32'h6f632720;
         'd3398: data <= 32'h6769666e;         'd3399: data <= 32'h41544f54;
         'd3400: data <= 32'h45485f4c;         'd3401: data <= 32'h535f5041;
         'd3402: data <= 32'h27455a49;         'd3403: data <= 32'h206e6920;
         'd3404: data <= 32'h65657246;         'd3405: data <= 32'h534f5452;
         'd3406: data <= 32'h666e6f43;         'd3407: data <= 32'h682e6769;
         'd3408: data <= 32'h00000a29;         'd3409: data <= 32'h65657246;
         'd3410: data <= 32'h534f5452;         'd3411: data <= 32'h5541465f;
         'd3412: data <= 32'h203a544c;         'd3413: data <= 32'h70704176;
         'd3414: data <= 32'h6163696c;         'd3415: data <= 32'h6e6f6974;
         'd3416: data <= 32'h63617453;         'd3417: data <= 32'h65764f6b;
         'd3418: data <= 32'h6f6c6672;         'd3419: data <= 32'h6f6f4877;
         'd3420: data <= 32'h00000a6b;         'd3421: data <= 32'hffffd200;
         'd3422: data <= 32'hffffd23c;         'd3423: data <= 32'hffffd23c;
         'd3424: data <= 32'hffffd23c;         'd3425: data <= 32'hffffd23c;
         'd3426: data <= 32'hffffd23c;         'd3427: data <= 32'hffffd23c;
         'd3428: data <= 32'hffffd23c;         'd3429: data <= 32'hffffd23c;
         'd3430: data <= 32'hffffd23c;         'd3431: data <= 32'hffffd23c;
         'd3432: data <= 32'hffffd188;         'd3433: data <= 32'hffffd1a0;
         'd3434: data <= 32'hffffd23c;         'd3435: data <= 32'hffffd23c;
         'd3436: data <= 32'hffffd23c;         'd3437: data <= 32'hffffd23c;
         'd3438: data <= 32'hffffd1a0;         'd3439: data <= 32'hffffd23c;
         'd3440: data <= 32'hffffd23c;         'd3441: data <= 32'hffffd23c;
         'd3442: data <= 32'hffffd23c;         'd3443: data <= 32'hffffd23c;
         'd3444: data <= 32'hffffd23c;         'd3445: data <= 32'hffffd200;
         'd3446: data <= 32'hffffd23c;         'd3447: data <= 32'hffffd23c;
         'd3448: data <= 32'hffffd170;         'd3449: data <= 32'hffffd23c;
         'd3450: data <= 32'hffffd1dc;         'd3451: data <= 32'hffffd23c;
         'd3452: data <= 32'hffffd23c;         'd3453: data <= 32'hffffd200;
         'd3454: data <= 32'h33323130;         'd3455: data <= 32'h37363534;
         'd3456: data <= 32'h62613938;         'd3457: data <= 32'h66656463;
         'd3458: data <= 32'h00000000;         'd3459: data <= 32'h33323130;
         'd3460: data <= 32'h37363534;         'd3461: data <= 32'h00003938;
         'd3462: data <= 32'h454c4449;         'd3463: data <= 32'h00000000;
         'd3464: data <= 32'hffffe6ec;         'd3465: data <= 32'hffffe768;
         'd3466: data <= 32'hffffe768;         'd3467: data <= 32'hffffe7d0;
         'd3468: data <= 32'hffffe7e0;         'd3469: data <= 32'hffffe81c;
         'd3470: data <= 32'hffffe768;         'd3471: data <= 32'hffffe768;
         'd3472: data <= 32'hffffe7d0;         'd3473: data <= 32'hffffe7e0;
         'd3474: data <= 32'h51726d54;         'd3475: data <= 32'h00000000;
         'd3476: data <= 32'h20726d54;         'd3477: data <= 32'h00637653;
         'd3478: data <= 32'h02020100;         'd3479: data <= 32'h03030303;
         'd3480: data <= 32'h04040404;         'd3481: data <= 32'h04040404;
         'd3482: data <= 32'h05050505;         'd3483: data <= 32'h05050505;
         'd3484: data <= 32'h05050505;         'd3485: data <= 32'h05050505;
         'd3486: data <= 32'h06060606;         'd3487: data <= 32'h06060606;
         'd3488: data <= 32'h06060606;         'd3489: data <= 32'h06060606;
         'd3490: data <= 32'h06060606;         'd3491: data <= 32'h06060606;
         'd3492: data <= 32'h06060606;         'd3493: data <= 32'h06060606;
         'd3494: data <= 32'h07070707;         'd3495: data <= 32'h07070707;
         'd3496: data <= 32'h07070707;         'd3497: data <= 32'h07070707;
         'd3498: data <= 32'h07070707;         'd3499: data <= 32'h07070707;
         'd3500: data <= 32'h07070707;         'd3501: data <= 32'h07070707;
         'd3502: data <= 32'h07070707;         'd3503: data <= 32'h07070707;
         'd3504: data <= 32'h07070707;         'd3505: data <= 32'h07070707;
         'd3506: data <= 32'h07070707;         'd3507: data <= 32'h07070707;
         'd3508: data <= 32'h07070707;         'd3509: data <= 32'h07070707;
         'd3510: data <= 32'h08080808;         'd3511: data <= 32'h08080808;
         'd3512: data <= 32'h08080808;         'd3513: data <= 32'h08080808;
         'd3514: data <= 32'h08080808;         'd3515: data <= 32'h08080808;
         'd3516: data <= 32'h08080808;         'd3517: data <= 32'h08080808;
         'd3518: data <= 32'h08080808;         'd3519: data <= 32'h08080808;
         'd3520: data <= 32'h08080808;         'd3521: data <= 32'h08080808;
         'd3522: data <= 32'h08080808;         'd3523: data <= 32'h08080808;
         'd3524: data <= 32'h08080808;         'd3525: data <= 32'h08080808;
         'd3526: data <= 32'h08080808;         'd3527: data <= 32'h08080808;
         'd3528: data <= 32'h08080808;         'd3529: data <= 32'h08080808;
         'd3530: data <= 32'h08080808;         'd3531: data <= 32'h08080808;
         'd3532: data <= 32'h08080808;         'd3533: data <= 32'h08080808;
         'd3534: data <= 32'h08080808;         'd3535: data <= 32'h08080808;
         'd3536: data <= 32'h08080808;         'd3537: data <= 32'h08080808;
         'd3538: data <= 32'h08080808;         'd3539: data <= 32'h08080808;
         'd3540: data <= 32'h08080808;         'd3541: data <= 32'h08080808;
         'd3542: data <= 32'h000186a0;         'd3543: data <= 32'h10001fd0;
         'd3544: data <= 32'h00000004;         'd3545: data <= 32'h10000010;
         'd3546: data <= 32'haaaaaaaa;         'd3547: data <= 32'h10000098;
         default: data <= '0;
         endcase
     end
 end
endmodule
